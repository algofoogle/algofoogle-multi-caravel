magic
tech gf180mcuD
magscale 1 5
timestamp 1702321337
<< metal2 >>
rect 5516 297836 5628 298500
rect 16548 297836 16660 298500
rect 27580 297836 27692 298500
rect 5502 297780 5628 297836
rect 16534 297780 16660 297836
rect 27566 297780 27692 297836
rect 38612 297836 38724 298500
rect 49644 297836 49756 298500
rect 60676 297836 60788 298500
rect 71708 297836 71820 298500
rect 82740 297836 82852 298500
rect 93772 297836 93884 298500
rect 104804 297836 104916 298500
rect 115836 297836 115948 298500
rect 126868 297836 126980 298500
rect 137900 297836 138012 298500
rect 148932 297836 149044 298500
rect 159964 297836 160076 298500
rect 38612 297780 38738 297836
rect 49644 297780 49770 297836
rect 60676 297780 60802 297836
rect 71708 297780 71834 297836
rect 82740 297780 82866 297836
rect 5502 156674 5530 297780
rect 16534 157234 16562 297780
rect 20398 295274 20426 295279
rect 20398 157794 20426 295246
rect 27566 295274 27594 297780
rect 27566 295241 27594 295246
rect 38710 295274 38738 297780
rect 49742 295330 49770 297780
rect 60774 295386 60802 297780
rect 71806 295442 71834 297780
rect 82838 295666 82866 297780
rect 93758 297780 93884 297836
rect 104790 297780 104916 297836
rect 115822 297780 115948 297836
rect 126854 297780 126980 297836
rect 137886 297780 138012 297836
rect 148918 297780 149044 297836
rect 159950 297780 160076 297836
rect 170996 297836 171108 298500
rect 182028 297836 182140 298500
rect 193060 297836 193172 298500
rect 204092 297836 204204 298500
rect 215124 297836 215236 298500
rect 226156 297836 226268 298500
rect 237188 297836 237300 298500
rect 248220 297836 248332 298500
rect 259252 297836 259364 298500
rect 170996 297780 171122 297836
rect 182028 297780 182154 297836
rect 193060 297780 193186 297836
rect 204092 297780 204218 297836
rect 82838 295633 82866 295638
rect 86926 295666 86954 295671
rect 71806 295409 71834 295414
rect 60774 295353 60802 295358
rect 86086 295386 86114 295391
rect 49742 295297 49770 295302
rect 38710 295241 38738 295246
rect 22918 168434 22946 170044
rect 22918 168401 22946 168406
rect 24262 161714 24290 170044
rect 25606 161770 25634 170044
rect 26950 166754 26978 170044
rect 26950 166721 26978 166726
rect 28294 161826 28322 170044
rect 29638 161882 29666 170044
rect 30982 164234 31010 170044
rect 30982 164201 31010 164206
rect 32326 162554 32354 170044
rect 32326 162521 32354 162526
rect 29638 161849 29666 161854
rect 28294 161793 28322 161798
rect 25606 161737 25634 161742
rect 24262 161681 24290 161686
rect 33670 161322 33698 170044
rect 33670 161289 33698 161294
rect 34062 168434 34090 168439
rect 34062 159964 34090 168406
rect 34734 161714 34762 161719
rect 34734 159964 34762 161686
rect 35014 161714 35042 170044
rect 36078 166754 36106 166759
rect 35014 161681 35042 161686
rect 35406 161770 35434 161775
rect 35406 159964 35434 161742
rect 36078 159964 36106 166726
rect 36358 162106 36386 170044
rect 36358 162073 36386 162078
rect 37422 161882 37450 161887
rect 36750 161826 36778 161831
rect 36750 159964 36778 161798
rect 37422 159964 37450 161854
rect 37702 161826 37730 170044
rect 37702 161793 37730 161798
rect 38094 164234 38122 164239
rect 38094 159964 38122 164206
rect 38766 162554 38794 162559
rect 38766 159964 38794 162526
rect 39046 161882 39074 170044
rect 39046 161849 39074 161854
rect 40110 161714 40138 161719
rect 39438 161322 39466 161327
rect 39438 159964 39466 161294
rect 40110 159964 40138 161686
rect 40390 161322 40418 170044
rect 41734 162162 41762 170044
rect 41734 162129 41762 162134
rect 40390 161289 40418 161294
rect 40782 162106 40810 162111
rect 40782 159964 40810 162078
rect 42126 161882 42154 161887
rect 41454 161826 41482 161831
rect 41454 159964 41482 161798
rect 42126 159964 42154 161854
rect 42798 161322 42826 161327
rect 42798 159964 42826 161294
rect 43078 161322 43106 170044
rect 43078 161289 43106 161294
rect 44142 162162 44170 162167
rect 44142 159964 44170 162134
rect 44422 162106 44450 170044
rect 45780 170030 46186 170058
rect 44422 162073 44450 162078
rect 45486 162106 45514 162111
rect 44814 161322 44842 161327
rect 44814 159964 44842 161294
rect 45486 159964 45514 162078
rect 46158 159964 46186 170030
rect 47110 168854 47138 170044
rect 47054 168826 47138 168854
rect 47054 167202 47082 168826
rect 48174 167258 48202 167263
rect 46830 167174 47082 167202
rect 47502 167202 47530 167207
rect 46830 159964 46858 167174
rect 47502 159964 47530 167174
rect 48174 159964 48202 167230
rect 48454 167202 48482 170044
rect 49798 167258 49826 170044
rect 49798 167225 49826 167230
rect 50190 167762 50218 167767
rect 48454 167169 48482 167174
rect 48846 167202 48874 167207
rect 48846 159964 48874 167174
rect 49518 163002 49546 163007
rect 49518 159964 49546 162974
rect 50190 159964 50218 167734
rect 50862 167706 50890 167711
rect 50862 159964 50890 167678
rect 51142 167202 51170 170044
rect 52206 167594 52234 167599
rect 51142 167169 51170 167174
rect 51534 167202 51562 167207
rect 51534 159964 51562 167174
rect 52206 159964 52234 167566
rect 52486 163002 52514 170044
rect 53830 167762 53858 170044
rect 53830 167729 53858 167734
rect 55174 167706 55202 170044
rect 55174 167673 55202 167678
rect 56518 167202 56546 170044
rect 57862 167594 57890 170044
rect 57862 167561 57890 167566
rect 56518 167169 56546 167174
rect 56910 167034 56938 167039
rect 53550 166922 53578 166927
rect 52486 162969 52514 162974
rect 52878 166754 52906 166759
rect 52878 159964 52906 166726
rect 53550 159964 53578 166894
rect 56238 161714 56266 161719
rect 56238 159964 56266 161686
rect 56910 159964 56938 167006
rect 57582 166978 57610 166983
rect 57582 159964 57610 166950
rect 58254 166866 58282 166871
rect 58254 159964 58282 166838
rect 58926 166810 58954 166815
rect 58926 159964 58954 166782
rect 59206 166754 59234 170044
rect 60270 168658 60298 168663
rect 59206 166721 59234 166726
rect 59598 166754 59626 166759
rect 59598 159964 59626 166726
rect 60270 159964 60298 168630
rect 60550 166922 60578 170044
rect 60550 166889 60578 166894
rect 60942 168602 60970 168607
rect 60942 159964 60970 168574
rect 61614 168434 61642 168439
rect 61614 159964 61642 168406
rect 61894 161714 61922 170044
rect 63238 167034 63266 170044
rect 63238 167001 63266 167006
rect 63406 168546 63434 168551
rect 61894 161681 61922 161686
rect 62286 162106 62314 162111
rect 62286 159964 62314 162078
rect 63406 162106 63434 168518
rect 63406 162073 63434 162078
rect 64414 168490 64442 168495
rect 62958 162050 62986 162055
rect 62958 159964 62986 162022
rect 64414 162050 64442 168462
rect 64582 166978 64610 170044
rect 64582 166945 64610 166950
rect 65926 166866 65954 170044
rect 65926 166833 65954 166838
rect 67270 166810 67298 170044
rect 67270 166777 67298 166782
rect 68614 166754 68642 170044
rect 69958 168658 69986 170044
rect 69958 168625 69986 168630
rect 71302 168602 71330 170044
rect 71302 168569 71330 168574
rect 72646 168434 72674 170044
rect 73990 168546 74018 170044
rect 73990 168513 74018 168518
rect 75334 168490 75362 170044
rect 75334 168457 75362 168462
rect 72646 168401 72674 168406
rect 68614 166721 68642 166726
rect 64414 162017 64442 162022
rect 70966 165074 70994 165079
rect 65646 161994 65674 161999
rect 63630 161938 63658 161943
rect 63630 159964 63658 161910
rect 64302 161882 64330 161887
rect 64302 159964 64330 161854
rect 64974 161826 65002 161831
rect 64974 159964 65002 161798
rect 65646 159964 65674 161966
rect 70966 161994 70994 165046
rect 70966 161961 70994 161966
rect 76678 161938 76706 170044
rect 76678 161905 76706 161910
rect 78022 161882 78050 170044
rect 78022 161849 78050 161854
rect 79366 161826 79394 170044
rect 80710 165074 80738 170044
rect 80710 165041 80738 165046
rect 79366 161793 79394 161798
rect 66318 161770 66346 161775
rect 66318 159964 66346 161742
rect 82054 161770 82082 170044
rect 82054 161737 82082 161742
rect 66990 161714 67018 161719
rect 66990 159964 67018 161686
rect 83398 161714 83426 170044
rect 86086 162106 86114 295358
rect 86086 162073 86114 162078
rect 86478 295274 86506 295279
rect 83398 161681 83426 161686
rect 86478 159964 86506 295246
rect 86926 161378 86954 295638
rect 86926 161345 86954 161350
rect 87038 295442 87066 295447
rect 87038 161322 87066 295414
rect 93646 295442 93674 295447
rect 87038 161289 87066 161294
rect 87150 295330 87178 295335
rect 87150 159964 87178 295302
rect 87822 162106 87850 162111
rect 87822 159964 87850 162078
rect 91854 162106 91882 162111
rect 89838 162050 89866 162055
rect 89166 161378 89194 161383
rect 88494 161322 88522 161327
rect 88494 159964 88522 161294
rect 89166 159964 89194 161350
rect 89838 159964 89866 162022
rect 90510 161826 90538 161831
rect 90510 159964 90538 161798
rect 91182 161714 91210 161719
rect 91182 159964 91210 161686
rect 91854 159964 91882 162078
rect 93646 162106 93674 295414
rect 93646 162073 93674 162078
rect 93758 162050 93786 297780
rect 95326 295554 95354 295559
rect 93758 162017 93786 162022
rect 93870 295274 93898 295279
rect 93198 161770 93226 161775
rect 92526 161322 92554 161327
rect 92526 159964 92554 161294
rect 93198 159964 93226 161742
rect 93870 159964 93898 295246
rect 95326 161826 95354 295526
rect 104790 295554 104818 297780
rect 104790 295521 104818 295526
rect 99526 295498 99554 295503
rect 95326 161793 95354 161798
rect 95438 295386 95466 295391
rect 95438 161322 95466 295358
rect 99526 161714 99554 295470
rect 115822 295498 115850 297780
rect 115822 295465 115850 295470
rect 126854 295442 126882 297780
rect 126854 295409 126882 295414
rect 137886 295386 137914 297780
rect 137886 295353 137914 295358
rect 99638 295330 99666 295335
rect 99638 161770 99666 295302
rect 148918 295330 148946 297780
rect 148918 295297 148946 295302
rect 159950 295274 159978 297780
rect 159950 295241 159978 295246
rect 171094 295274 171122 297780
rect 182126 295330 182154 297780
rect 193158 295386 193186 297780
rect 204190 295442 204218 297780
rect 204190 295409 204218 295414
rect 215110 297780 215236 297836
rect 226142 297780 226268 297836
rect 237174 297780 237300 297836
rect 248206 297780 248332 297836
rect 259238 297780 259364 297836
rect 269710 297822 270242 297850
rect 270284 297836 270396 298500
rect 281316 297836 281428 298500
rect 292348 297836 292460 298500
rect 193158 295353 193186 295358
rect 182126 295297 182154 295302
rect 208726 295330 208754 295335
rect 171094 295241 171122 295246
rect 102606 167314 102634 167319
rect 99638 161737 99666 161742
rect 101934 167202 101962 167207
rect 99526 161681 99554 161686
rect 95438 161289 95466 161294
rect 101934 159964 101962 167174
rect 102606 159964 102634 167286
rect 102942 167202 102970 170044
rect 102942 167169 102970 167174
rect 103278 167370 103306 167375
rect 103278 159964 103306 167342
rect 104286 167314 104314 170044
rect 104286 167281 104314 167286
rect 105294 168042 105322 168047
rect 104622 163786 104650 163791
rect 103950 163450 103978 163455
rect 103950 159964 103978 163422
rect 104622 159964 104650 163758
rect 105294 159964 105322 168014
rect 105630 167370 105658 170044
rect 106638 167930 106666 167935
rect 105630 167337 105658 167342
rect 105966 167370 105994 167375
rect 105966 159964 105994 167342
rect 106638 159964 106666 167902
rect 106974 163450 107002 170044
rect 106974 163417 107002 163422
rect 107310 167874 107338 167879
rect 107310 159964 107338 167846
rect 107982 167818 108010 167823
rect 107982 159964 108010 167790
rect 108318 163786 108346 170044
rect 109662 168042 109690 170044
rect 109662 168009 109690 168014
rect 108318 163753 108346 163758
rect 108654 167762 108682 167767
rect 108654 159964 108682 167734
rect 109326 167706 109354 167711
rect 109326 159964 109354 167678
rect 109998 167650 110026 167655
rect 109998 159964 110026 167622
rect 111006 167370 111034 170044
rect 112350 167930 112378 170044
rect 112350 167897 112378 167902
rect 113694 167874 113722 170044
rect 113694 167841 113722 167846
rect 114702 168658 114730 168663
rect 111006 167337 111034 167342
rect 112014 167594 112042 167599
rect 110670 161882 110698 161887
rect 110670 159964 110698 161854
rect 112014 159964 112042 167566
rect 112686 162554 112714 162559
rect 112686 159964 112714 162526
rect 113358 161826 113386 161831
rect 113358 159964 113386 161798
rect 114030 161770 114058 161775
rect 114030 159964 114058 161742
rect 114702 159964 114730 168630
rect 115038 167818 115066 170044
rect 115038 167785 115066 167790
rect 116046 168602 116074 168607
rect 115374 161714 115402 161719
rect 115374 159964 115402 161686
rect 116046 159964 116074 168574
rect 116382 167762 116410 170044
rect 116382 167729 116410 167734
rect 116718 168546 116746 168551
rect 116718 159964 116746 168518
rect 117390 168490 117418 168495
rect 116774 163786 116802 163791
rect 116774 161882 116802 163758
rect 116774 161849 116802 161854
rect 117390 159964 117418 168462
rect 117726 167706 117754 170044
rect 117726 167673 117754 167678
rect 118062 168434 118090 168439
rect 118062 159964 118090 168406
rect 119070 167650 119098 170044
rect 119070 167617 119098 167622
rect 120414 163786 120442 170044
rect 121758 167594 121786 170044
rect 121758 167561 121786 167566
rect 120414 163753 120442 163758
rect 120078 163450 120106 163455
rect 118734 162106 118762 162111
rect 118734 159964 118762 162078
rect 119406 162050 119434 162055
rect 119406 159964 119434 162022
rect 120078 159964 120106 163422
rect 121422 163394 121450 163399
rect 120750 161938 120778 161943
rect 120750 159964 120778 161910
rect 121422 159964 121450 163366
rect 123102 162554 123130 170044
rect 123102 162521 123130 162526
rect 124110 161994 124138 161999
rect 124110 159964 124138 161966
rect 124446 161826 124474 170044
rect 125566 168714 125594 168719
rect 125566 162106 125594 168686
rect 125566 162073 125594 162078
rect 124446 161793 124474 161798
rect 125454 161882 125482 161887
rect 124782 161658 124810 161663
rect 124782 159964 124810 161630
rect 125454 159964 125482 161854
rect 125790 161770 125818 170044
rect 127134 168658 127162 170044
rect 127134 168625 127162 168630
rect 127470 162666 127498 162671
rect 125790 161737 125818 161742
rect 126126 162554 126154 162559
rect 126126 159964 126154 162526
rect 126798 161826 126826 161831
rect 126798 159964 126826 161798
rect 127470 159964 127498 162638
rect 128142 161770 128170 161775
rect 128142 159964 128170 161742
rect 128478 161714 128506 170044
rect 129822 168602 129850 170044
rect 129822 168569 129850 168574
rect 129934 168658 129962 168663
rect 128478 161681 128506 161686
rect 128814 162610 128842 162615
rect 128814 159964 128842 162582
rect 129486 161714 129514 161719
rect 129486 159964 129514 161686
rect 129934 161658 129962 168630
rect 131166 168546 131194 170044
rect 131166 168513 131194 168518
rect 131614 168602 131642 168607
rect 130830 162890 130858 162895
rect 129934 161625 129962 161630
rect 130158 162162 130186 162167
rect 130158 159964 130186 162134
rect 130830 159964 130858 162862
rect 131502 162834 131530 162839
rect 131502 159964 131530 162806
rect 131614 162554 131642 168574
rect 132286 168546 132314 168551
rect 131614 162521 131642 162526
rect 132174 162778 132202 162783
rect 132174 159964 132202 162750
rect 132286 162666 132314 168518
rect 132510 168490 132538 170044
rect 132510 168457 132538 168462
rect 133854 168434 133882 170044
rect 135198 168714 135226 170044
rect 135198 168681 135226 168686
rect 133854 168401 133882 168406
rect 133966 168490 133994 168495
rect 132286 162633 132314 162638
rect 132846 162722 132874 162727
rect 132846 159964 132874 162694
rect 133518 162666 133546 162671
rect 133518 159964 133546 162638
rect 133966 162610 133994 168462
rect 134974 168434 135002 168439
rect 133966 162577 133994 162582
rect 134190 162610 134218 162615
rect 134190 159964 134218 162582
rect 134862 162554 134890 162559
rect 134862 159964 134890 162526
rect 134974 162162 135002 168406
rect 134974 162129 135002 162134
rect 136542 162050 136570 170044
rect 137886 163450 137914 170044
rect 137886 163417 137914 163422
rect 136542 162017 136570 162022
rect 139230 161938 139258 170044
rect 140574 163394 140602 170044
rect 140574 163361 140602 163366
rect 141918 161994 141946 170044
rect 143262 168658 143290 170044
rect 143262 168625 143290 168630
rect 141918 161961 141946 161966
rect 139230 161905 139258 161910
rect 144606 161882 144634 170044
rect 145950 168602 145978 170044
rect 145950 168569 145978 168574
rect 144606 161849 144634 161854
rect 147294 161826 147322 170044
rect 148638 168546 148666 170044
rect 148638 168513 148666 168518
rect 147294 161793 147322 161798
rect 149982 161770 150010 170044
rect 151326 168490 151354 170044
rect 151326 168457 151354 168462
rect 149982 161737 150010 161742
rect 152670 161714 152698 170044
rect 154014 168434 154042 170044
rect 154014 168401 154042 168406
rect 155358 162890 155386 170044
rect 155358 162857 155386 162862
rect 156702 162834 156730 170044
rect 156702 162801 156730 162806
rect 158046 162778 158074 170044
rect 158046 162745 158074 162750
rect 159390 162722 159418 170044
rect 159390 162689 159418 162694
rect 160734 162666 160762 170044
rect 160734 162633 160762 162638
rect 162078 162610 162106 170044
rect 162078 162577 162106 162582
rect 163422 162554 163450 170044
rect 180558 168602 180586 168607
rect 179886 168546 179914 168551
rect 179214 168490 179242 168495
rect 175854 168434 175882 168439
rect 163422 162521 163450 162526
rect 174510 167594 174538 167599
rect 152670 161681 152698 161686
rect 174510 159964 174538 167566
rect 175182 165914 175210 165919
rect 175182 159964 175210 165886
rect 175854 159964 175882 168406
rect 179214 159964 179242 168462
rect 179886 159964 179914 168518
rect 180558 159964 180586 168574
rect 181006 167594 181034 170044
rect 181006 167561 181034 167566
rect 181230 167258 181258 167263
rect 181230 159964 181258 167230
rect 181566 165914 181594 170044
rect 181566 165881 181594 165886
rect 181902 167202 181930 167207
rect 181902 159964 181930 167174
rect 182126 164626 182154 170044
rect 182126 164593 182154 164598
rect 182574 164626 182602 164631
rect 182574 159964 182602 164598
rect 182686 164626 182714 170044
rect 183260 170030 183722 170058
rect 182686 164593 182714 164598
rect 183246 164626 183274 164631
rect 183246 159964 183274 164598
rect 183694 159978 183722 170030
rect 183806 167258 183834 170044
rect 183806 167225 183834 167230
rect 184366 167202 184394 170044
rect 184814 170030 184940 170058
rect 185262 170030 185500 170058
rect 185934 170030 186060 170058
rect 184814 167202 184842 170030
rect 184366 167169 184394 167174
rect 184590 167174 184842 167202
rect 183694 159950 183932 159978
rect 184590 159964 184618 167174
rect 185262 159964 185290 170030
rect 185934 159964 185962 170030
rect 186606 159964 186634 170044
rect 187180 170030 187306 170058
rect 187278 159964 187306 170030
rect 187726 168434 187754 170044
rect 188286 168546 188314 170044
rect 188846 168602 188874 170044
rect 188846 168569 188874 168574
rect 188286 168513 188314 168518
rect 187726 168401 187754 168406
rect 187950 167258 187978 167263
rect 187950 159964 187978 167230
rect 189406 167258 189434 170044
rect 189406 167225 189434 167230
rect 188622 167202 188650 167207
rect 188622 159964 188650 167174
rect 189966 167202 189994 170044
rect 190526 168490 190554 170044
rect 190526 168457 190554 168462
rect 189966 167169 189994 167174
rect 191086 162050 191114 170044
rect 191646 168658 191674 170044
rect 191646 168625 191674 168630
rect 191086 162017 191114 162022
rect 192206 161994 192234 170044
rect 192206 161961 192234 161966
rect 192766 161938 192794 170044
rect 192766 161905 192794 161910
rect 193326 161882 193354 170044
rect 193886 168546 193914 170044
rect 193886 168513 193914 168518
rect 193326 161849 193354 161854
rect 194446 161826 194474 170044
rect 195006 168490 195034 170044
rect 195006 168457 195034 168462
rect 194446 161793 194474 161798
rect 195566 161770 195594 170044
rect 196126 168434 196154 170044
rect 196126 168401 196154 168406
rect 195566 161737 195594 161742
rect 196686 161714 196714 170044
rect 197246 168602 197274 170044
rect 197246 168569 197274 168574
rect 197806 162666 197834 170044
rect 198366 168714 198394 170044
rect 198366 168681 198394 168686
rect 197806 162633 197834 162638
rect 198926 162554 198954 170044
rect 199486 168770 199514 170044
rect 199486 168737 199514 168742
rect 198926 162521 198954 162526
rect 200046 162498 200074 170044
rect 200046 162465 200074 162470
rect 200606 162442 200634 170044
rect 201166 162890 201194 170044
rect 201166 162857 201194 162862
rect 201726 162834 201754 170044
rect 201726 162801 201754 162806
rect 202062 168658 202090 168663
rect 200606 162409 200634 162414
rect 201166 162666 201194 162671
rect 201166 162106 201194 162638
rect 201166 162073 201194 162078
rect 196686 161681 196714 161686
rect 201390 162050 201418 162055
rect 201390 159964 201418 162022
rect 202062 159964 202090 168630
rect 202286 162778 202314 170044
rect 202286 162745 202314 162750
rect 202846 162722 202874 170044
rect 202846 162689 202874 162694
rect 203406 162666 203434 170044
rect 203406 162633 203434 162638
rect 202454 162554 202482 162559
rect 202454 162050 202482 162526
rect 203966 162554 203994 170044
rect 205534 168770 205562 168775
rect 203966 162521 203994 162526
rect 204750 168546 204778 168551
rect 202454 162017 202482 162022
rect 203294 162498 203322 162503
rect 202734 161994 202762 161999
rect 202734 159964 202762 161966
rect 203294 161994 203322 162470
rect 203294 161961 203322 161966
rect 203518 162442 203546 162447
rect 203406 161938 203434 161943
rect 203406 159964 203434 161910
rect 203518 161938 203546 162414
rect 203518 161905 203546 161910
rect 204078 161882 204106 161887
rect 204078 159964 204106 161854
rect 204750 159964 204778 168518
rect 205422 161826 205450 161831
rect 205422 159964 205450 161798
rect 205534 161826 205562 168742
rect 207046 168714 207074 168719
rect 205534 161793 205562 161798
rect 206094 168490 206122 168495
rect 206094 159964 206122 168462
rect 207046 162974 207074 168686
rect 207886 168602 207914 168607
rect 207438 168434 207466 168439
rect 207046 162946 207186 162974
rect 207158 162050 207186 162946
rect 207158 162017 207186 162022
rect 206766 161770 206794 161775
rect 206766 159964 206794 161742
rect 207438 159964 207466 168406
rect 207886 161322 207914 168574
rect 208726 162610 208754 295302
rect 215110 166754 215138 297780
rect 216398 295442 216426 295447
rect 215110 166721 215138 166726
rect 216286 295386 216314 295391
rect 208726 162577 208754 162582
rect 213486 162890 213514 162895
rect 209454 162106 209482 162111
rect 207886 161289 207914 161294
rect 208110 161714 208138 161719
rect 208110 159964 208138 161686
rect 208782 161322 208810 161327
rect 208782 159964 208810 161294
rect 209454 159964 209482 162078
rect 210126 162050 210154 162055
rect 210126 159964 210154 162022
rect 212142 161994 212170 161999
rect 211470 161826 211498 161831
rect 210798 161770 210826 161775
rect 210798 159964 210826 161742
rect 211470 159964 211498 161798
rect 212142 159964 212170 161966
rect 212814 161938 212842 161943
rect 212814 159964 212842 161910
rect 213486 159964 213514 162862
rect 214158 162834 214186 162839
rect 214158 159964 214186 162806
rect 214830 162778 214858 162783
rect 214830 159964 214858 162750
rect 215502 162722 215530 162727
rect 215502 159964 215530 162694
rect 216174 162666 216202 162671
rect 216174 159964 216202 162638
rect 216286 161770 216314 295358
rect 216286 161737 216314 161742
rect 216398 161714 216426 295414
rect 225582 295330 225610 295335
rect 216398 161681 216426 161686
rect 216510 295274 216538 295279
rect 216510 161322 216538 295246
rect 224686 295106 224714 295111
rect 223566 166754 223594 166759
rect 221550 162610 221578 162615
rect 216510 161289 216538 161294
rect 216846 162554 216874 162559
rect 216846 159964 216874 162526
rect 220878 161322 220906 161327
rect 220878 159964 220906 161294
rect 221550 159964 221578 162582
rect 222222 161770 222250 161775
rect 222222 159964 222250 161742
rect 222894 161714 222922 161719
rect 222894 159964 222922 161686
rect 223566 159964 223594 166726
rect 224238 161322 224266 161327
rect 224238 159964 224266 161294
rect 224686 161322 224714 295078
rect 224686 161289 224714 161294
rect 224910 161322 224938 161327
rect 224910 159964 224938 161294
rect 225582 159964 225610 295302
rect 226142 295106 226170 297780
rect 227206 295386 227234 295391
rect 226142 295073 226170 295078
rect 226254 295274 226282 295279
rect 226254 159964 226282 295246
rect 227206 161322 227234 295358
rect 237174 295386 237202 297780
rect 237174 295353 237202 295358
rect 248206 295330 248234 297780
rect 248206 295297 248234 295302
rect 259238 295274 259266 297780
rect 259238 295241 259266 295246
rect 235662 166306 235690 166311
rect 232974 166250 233002 166255
rect 232302 165970 232330 165975
rect 227206 161289 227234 161294
rect 230286 165914 230314 165919
rect 230286 159964 230314 165886
rect 230958 161714 230986 161719
rect 230958 159964 230986 161686
rect 232302 159964 232330 165942
rect 232974 159964 233002 166222
rect 234990 166194 235018 166199
rect 233646 165858 233674 165863
rect 233646 159964 233674 165830
rect 234318 165802 234346 165807
rect 234318 159964 234346 165774
rect 234990 159964 235018 166166
rect 235662 159964 235690 166278
rect 235886 165914 235914 170044
rect 235886 165881 235914 165886
rect 236334 167762 236362 167767
rect 236334 159964 236362 167734
rect 236558 161714 236586 170044
rect 236558 161681 236586 161686
rect 237006 167650 237034 167655
rect 237006 159964 237034 167622
rect 237230 165970 237258 170044
rect 237230 165937 237258 165942
rect 237678 167594 237706 167599
rect 237678 159964 237706 167566
rect 237902 166250 237930 170044
rect 237902 166217 237930 166222
rect 238350 167706 238378 167711
rect 238350 159964 238378 167678
rect 238574 165858 238602 170044
rect 238574 165825 238602 165830
rect 239022 167986 239050 167991
rect 239022 159964 239050 167958
rect 239246 165802 239274 170044
rect 239246 165769 239274 165774
rect 239694 167202 239722 167207
rect 239694 159964 239722 167174
rect 239918 166194 239946 170044
rect 239918 166161 239946 166166
rect 240366 167930 240394 167935
rect 240366 159964 240394 167902
rect 240590 166306 240618 170044
rect 240590 166273 240618 166278
rect 241038 167874 241066 167879
rect 241038 159964 241066 167846
rect 241262 167762 241290 170044
rect 241262 167729 241290 167734
rect 241934 167650 241962 170044
rect 241934 167617 241962 167622
rect 242606 167594 242634 170044
rect 243278 167706 243306 170044
rect 243950 167986 243978 170044
rect 243950 167953 243978 167958
rect 243278 167673 243306 167678
rect 242606 167561 242634 167566
rect 244622 167202 244650 170044
rect 245294 167930 245322 170044
rect 245294 167897 245322 167902
rect 245966 167874 245994 170044
rect 245966 167841 245994 167846
rect 244622 167169 244650 167174
rect 246638 164234 246666 170044
rect 247310 164346 247338 170044
rect 247982 166026 248010 170044
rect 247982 165993 248010 165998
rect 248654 165914 248682 170044
rect 248654 165881 248682 165886
rect 247310 164313 247338 164318
rect 246638 164201 246666 164206
rect 249326 163450 249354 170044
rect 249998 164290 250026 170044
rect 249998 164257 250026 164262
rect 249326 163417 249354 163422
rect 250670 163394 250698 170044
rect 251342 165970 251370 170044
rect 251342 165937 251370 165942
rect 250670 163361 250698 163366
rect 252014 162554 252042 170044
rect 252686 162610 252714 170044
rect 253358 165074 253386 170044
rect 253358 165041 253386 165046
rect 253806 164346 253834 164351
rect 252686 162577 252714 162582
rect 253134 164234 253162 164239
rect 252014 162521 252042 162526
rect 253134 159964 253162 164206
rect 253806 159964 253834 164318
rect 254030 163506 254058 170044
rect 254702 168434 254730 170044
rect 254702 168401 254730 168406
rect 261198 168434 261226 168439
rect 254030 163473 254058 163478
rect 254478 166026 254506 166031
rect 254478 159964 254506 165998
rect 257838 165970 257866 165975
rect 255150 165914 255178 165919
rect 255150 159964 255178 165886
rect 256494 164290 256522 164295
rect 255822 163450 255850 163455
rect 255822 159964 255850 163422
rect 256494 159964 256522 164262
rect 257166 163394 257194 163399
rect 257166 159964 257194 163366
rect 257838 159964 257866 165942
rect 259854 165074 259882 165079
rect 259182 162610 259210 162615
rect 258510 162554 258538 162559
rect 258510 159964 258538 162526
rect 259182 159964 259210 162582
rect 259854 159964 259882 165046
rect 260526 163506 260554 163511
rect 260526 159964 260554 163478
rect 261198 159964 261226 168406
rect 269710 159362 269738 297822
rect 270214 297738 270242 297822
rect 270270 297780 270396 297836
rect 281302 297780 281428 297836
rect 292334 297780 292460 297836
rect 270270 297738 270298 297780
rect 270214 297710 270298 297738
rect 269710 159329 269738 159334
rect 273406 295274 273434 295279
rect 273406 158578 273434 295246
rect 281302 295274 281330 297780
rect 281302 295241 281330 295246
rect 273406 158545 273434 158550
rect 292334 158130 292362 297780
rect 292334 158097 292362 158102
rect 20398 157761 20426 157766
rect 16534 157201 16562 157206
rect 5502 156641 5530 156646
rect 277606 137522 277634 137527
rect 275422 135674 275450 135679
rect 272118 135282 272146 135287
rect 33950 129066 33978 129071
rect 16814 129010 16842 129015
rect 16814 104972 16842 128982
rect 24430 107114 24458 107119
rect 22526 106386 22554 106391
rect 18718 106330 18746 106335
rect 18718 104972 18746 106302
rect 20622 106274 20650 106279
rect 20622 104972 20650 106246
rect 22526 104972 22554 106358
rect 24430 104972 24458 107086
rect 30142 106610 30170 106615
rect 28238 106498 28266 106503
rect 26334 106442 26362 106447
rect 26334 104972 26362 106414
rect 28238 104972 28266 106470
rect 30142 104972 30170 106582
rect 32046 106554 32074 106559
rect 32046 104972 32074 106526
rect 33950 104972 33978 129038
rect 35070 129010 35098 130060
rect 35070 128977 35098 128982
rect 34846 128954 34874 128959
rect 34846 106330 34874 128926
rect 34846 106297 34874 106302
rect 35854 107170 35882 107175
rect 35854 104972 35882 107142
rect 37086 106274 37114 130060
rect 37366 129010 37394 129015
rect 37366 106610 37394 128982
rect 37366 106577 37394 106582
rect 37758 106386 37786 130060
rect 39102 106442 39130 130060
rect 39102 106409 39130 106414
rect 39662 106610 39690 106615
rect 37758 106353 37786 106358
rect 37086 106241 37114 106246
rect 37758 106274 37786 106279
rect 37758 104972 37786 106246
rect 39662 104972 39690 106582
rect 39774 106498 39802 130060
rect 41118 106554 41146 130060
rect 41790 129066 41818 130060
rect 41790 129033 41818 129038
rect 41118 106521 41146 106526
rect 41566 107226 41594 107231
rect 39774 106465 39802 106470
rect 41566 104972 41594 107198
rect 43134 106274 43162 130060
rect 43134 106241 43162 106246
rect 43470 106666 43498 106671
rect 43470 104972 43498 106638
rect 43806 106610 43834 130060
rect 45150 106666 45178 130060
rect 45150 106633 45178 106638
rect 45374 130046 45836 130074
rect 43806 106577 43834 106582
rect 45374 104972 45402 130046
rect 47166 106666 47194 130060
rect 47838 128898 47866 130060
rect 47838 128865 47866 128870
rect 48286 128898 48314 128903
rect 47166 106633 47194 106638
rect 47278 107282 47306 107287
rect 47278 104972 47306 107254
rect 48286 106610 48314 128870
rect 49182 128898 49210 130060
rect 49182 128865 49210 128870
rect 48286 106577 48314 106582
rect 49182 106666 49210 106671
rect 49182 104972 49210 106638
rect 49854 106330 49882 130060
rect 49966 128898 49994 128903
rect 49966 106386 49994 128870
rect 51198 128562 51226 130060
rect 51198 128529 51226 128534
rect 51646 128562 51674 128567
rect 49966 106353 49994 106358
rect 51086 106610 51114 106615
rect 49854 106297 49882 106302
rect 51086 104972 51114 106582
rect 51646 106274 51674 128534
rect 51870 106610 51898 130060
rect 51870 106577 51898 106582
rect 52990 107338 53018 107343
rect 51646 106241 51674 106246
rect 52990 104972 53018 107310
rect 53214 106442 53242 130060
rect 53886 129066 53914 130060
rect 53886 129033 53914 129038
rect 55230 106554 55258 130060
rect 55902 129122 55930 130060
rect 55902 129089 55930 129094
rect 57246 107394 57274 130060
rect 57246 107361 57274 107366
rect 55230 106521 55258 106526
rect 57918 106498 57946 130060
rect 57918 106465 57946 106470
rect 58702 107450 58730 107455
rect 53214 106409 53242 106414
rect 54894 106386 54922 106391
rect 54894 104972 54922 106358
rect 56798 106330 56826 106335
rect 56798 104972 56826 106302
rect 58702 104972 58730 107422
rect 59262 106386 59290 130060
rect 59262 106353 59290 106358
rect 59934 106330 59962 130060
rect 59934 106297 59962 106302
rect 60606 106274 60634 106279
rect 60606 104972 60634 106246
rect 61278 106274 61306 130060
rect 61950 129234 61978 130060
rect 61950 129201 61978 129206
rect 66990 129234 67018 129239
rect 66766 129178 66794 129183
rect 64414 106666 64442 106671
rect 61278 106241 61306 106246
rect 62510 106610 62538 106615
rect 62510 104972 62538 106582
rect 64414 104972 64442 106638
rect 66766 106666 66794 129150
rect 66766 106633 66794 106638
rect 66878 129066 66906 129071
rect 66878 106666 66906 129038
rect 66878 106633 66906 106638
rect 66318 106442 66346 106447
rect 66318 104972 66346 106414
rect 66990 106442 67018 129206
rect 68446 129122 68474 129127
rect 66990 106409 67018 106414
rect 68222 106666 68250 106671
rect 68222 104972 68250 106638
rect 68446 106610 68474 129094
rect 68446 106577 68474 106582
rect 70126 129066 70154 129071
rect 70126 104972 70154 129038
rect 70686 128954 70714 130060
rect 70686 128921 70714 128926
rect 71358 107114 71386 130060
rect 72030 129010 72058 130060
rect 72030 128977 72058 128982
rect 72702 107170 72730 130060
rect 73374 107226 73402 130060
rect 74046 107282 74074 130060
rect 74718 107338 74746 130060
rect 75390 107450 75418 130060
rect 76062 129178 76090 130060
rect 76062 129145 76090 129150
rect 76734 129066 76762 130060
rect 76734 129033 76762 129038
rect 75390 107417 75418 107422
rect 75838 128898 75866 128903
rect 74718 107305 74746 107310
rect 74046 107249 74074 107254
rect 73374 107193 73402 107198
rect 72702 107137 72730 107142
rect 71358 107081 71386 107086
rect 73934 106610 73962 106615
rect 72030 106554 72058 106559
rect 72030 104972 72058 106526
rect 73934 104972 73962 106582
rect 75838 104972 75866 128870
rect 77406 128898 77434 130060
rect 77406 128865 77434 128870
rect 77742 107394 77770 107399
rect 77742 104972 77770 107366
rect 78078 106666 78106 130060
rect 78078 106633 78106 106638
rect 78750 106554 78778 130060
rect 82782 127274 82810 130060
rect 82782 127241 82810 127246
rect 83454 126602 83482 130060
rect 84798 127330 84826 130060
rect 84798 127297 84826 127302
rect 83454 126569 83482 126574
rect 85470 126434 85498 130060
rect 86142 128954 86170 130060
rect 86142 128921 86170 128926
rect 86814 127386 86842 130060
rect 86814 127353 86842 127358
rect 87486 126490 87514 130060
rect 88158 126546 88186 130060
rect 88830 127442 88858 130060
rect 89502 128114 89530 130060
rect 90174 129010 90202 130060
rect 90174 128977 90202 128982
rect 89502 128081 89530 128086
rect 88830 127409 88858 127414
rect 90846 126770 90874 130060
rect 91518 129234 91546 130060
rect 91518 129201 91546 129206
rect 90846 126737 90874 126742
rect 92190 126658 92218 130060
rect 92862 127498 92890 130060
rect 93534 128170 93562 130060
rect 94206 129066 94234 130060
rect 94206 129033 94234 129038
rect 93534 128137 93562 128142
rect 92862 127465 92890 127470
rect 92190 126625 92218 126630
rect 88158 126513 88186 126518
rect 87486 126457 87514 126462
rect 85470 126401 85498 126406
rect 94878 126378 94906 130060
rect 95550 129290 95578 130060
rect 95550 129257 95578 129262
rect 96222 126714 96250 130060
rect 96894 129178 96922 130060
rect 97566 129346 97594 130060
rect 97566 129313 97594 129318
rect 96894 129145 96922 129150
rect 98238 129122 98266 130060
rect 98238 129089 98266 129094
rect 98910 128394 98938 130060
rect 98910 128361 98938 128366
rect 99134 129234 99162 129239
rect 99134 127554 99162 129206
rect 99582 128226 99610 130060
rect 99582 128193 99610 128198
rect 99134 127521 99162 127526
rect 100254 126826 100282 130060
rect 100926 129234 100954 130060
rect 100926 129201 100954 129206
rect 101598 128282 101626 130060
rect 101598 128249 101626 128254
rect 100254 126793 100282 126798
rect 102046 127274 102074 127279
rect 96222 126681 96250 126686
rect 94878 126345 94906 126350
rect 102046 124964 102074 127246
rect 102270 127274 102298 130060
rect 102886 129346 102914 129351
rect 102438 129290 102466 129295
rect 102438 127610 102466 129262
rect 102886 127666 102914 129318
rect 102886 127633 102914 127638
rect 102438 127577 102466 127582
rect 102270 127241 102298 127246
rect 102494 127330 102522 127335
rect 102270 126602 102298 126607
rect 102270 124964 102298 126574
rect 102494 124964 102522 127302
rect 102942 127218 102970 130060
rect 102942 127185 102970 127190
rect 103166 127386 103194 127391
rect 103166 124964 103194 127358
rect 103614 126602 103642 130060
rect 103614 126569 103642 126574
rect 103838 127442 103866 127447
rect 103838 124964 103866 127414
rect 104286 126322 104314 130060
rect 104958 126882 104986 130060
rect 104958 126849 104986 126854
rect 105182 127498 105210 127503
rect 104286 126289 104314 126294
rect 104510 126770 104538 126775
rect 104510 124964 104538 126742
rect 105182 124964 105210 127470
rect 105630 127330 105658 130060
rect 106302 128338 106330 130060
rect 106302 128305 106330 128310
rect 106526 129178 106554 129183
rect 105630 127297 105658 127302
rect 105854 126378 105882 126383
rect 105854 124964 105882 126350
rect 106526 124964 106554 129150
rect 106806 129010 106834 129015
rect 106806 128506 106834 128982
rect 106806 128473 106834 128478
rect 106974 126154 107002 130060
rect 106974 126121 107002 126126
rect 107198 128394 107226 128399
rect 107198 124964 107226 128366
rect 107646 127386 107674 130060
rect 107646 127353 107674 127358
rect 107870 129234 107898 129239
rect 107870 124964 107898 129206
rect 108150 128954 108178 128959
rect 108094 126434 108122 126439
rect 108094 124964 108122 126406
rect 108150 124978 108178 128926
rect 108318 127442 108346 130060
rect 108318 127409 108346 127414
rect 108542 127218 108570 127223
rect 108150 124950 108332 124978
rect 108542 124964 108570 127190
rect 108990 126770 109018 130060
rect 108990 126737 109018 126742
rect 109046 129066 109074 129071
rect 108990 126546 109018 126551
rect 108766 126490 108794 126495
rect 108766 124964 108794 126462
rect 108990 124964 109018 126518
rect 109046 126490 109074 129038
rect 109494 128506 109522 128511
rect 109438 128114 109466 128119
rect 109046 126457 109074 126462
rect 109214 126882 109242 126887
rect 109214 124964 109242 126854
rect 109438 124964 109466 128086
rect 109494 124978 109522 128478
rect 109662 127498 109690 130060
rect 109662 127465 109690 127470
rect 110054 129122 110082 129127
rect 109886 126154 109914 126159
rect 109494 124950 109676 124978
rect 109886 124964 109914 126126
rect 110054 126154 110082 129094
rect 110334 127694 110362 130060
rect 111020 130046 111258 130074
rect 110782 128170 110810 128175
rect 110334 127666 110418 127694
rect 110054 126121 110082 126126
rect 110110 127554 110138 127559
rect 110110 124964 110138 127526
rect 110334 126658 110362 126663
rect 110334 124964 110362 126630
rect 110390 126434 110418 127666
rect 110390 126401 110418 126406
rect 110558 126770 110586 126775
rect 110558 124964 110586 126742
rect 110782 124964 110810 128142
rect 111006 126490 111034 126495
rect 111006 124964 111034 126462
rect 111230 124964 111258 130046
rect 111678 128170 111706 130060
rect 112350 128674 112378 130060
rect 112350 128641 112378 128646
rect 112574 128898 112602 128903
rect 111678 128137 111706 128142
rect 112126 127666 112154 127671
rect 111454 127610 111482 127615
rect 111454 124964 111482 127582
rect 111902 126882 111930 126887
rect 111678 126378 111706 126383
rect 111678 124964 111706 126350
rect 111902 124964 111930 126854
rect 112126 124964 112154 127638
rect 112350 126154 112378 126159
rect 112350 124964 112378 126126
rect 112574 124964 112602 128870
rect 112798 128226 112826 128231
rect 112798 124964 112826 128198
rect 113022 126882 113050 130060
rect 113708 130046 113778 130074
rect 113022 126849 113050 126854
rect 113246 128618 113274 128623
rect 112854 126826 112882 126831
rect 112854 124978 112882 126798
rect 112854 124950 113036 124978
rect 113246 124964 113274 128590
rect 113470 128282 113498 128287
rect 113470 124964 113498 128254
rect 113694 127274 113722 127279
rect 113694 124964 113722 127246
rect 113750 126826 113778 130046
rect 113750 126793 113778 126798
rect 114142 126602 114170 126607
rect 113918 126490 113946 126495
rect 113918 124964 113946 126462
rect 114142 124964 114170 126574
rect 114366 126602 114394 130060
rect 114366 126569 114394 126574
rect 114590 129066 114618 129071
rect 114366 126322 114394 126327
rect 114366 124964 114394 126294
rect 114590 124964 114618 129038
rect 115038 128898 115066 130060
rect 115038 128865 115066 128870
rect 115262 129010 115290 129015
rect 115038 128338 115066 128343
rect 114814 127330 114842 127335
rect 114814 124964 114842 127302
rect 115038 124964 115066 128310
rect 115262 124964 115290 128982
rect 115542 127442 115570 127447
rect 115486 127386 115514 127391
rect 115486 124964 115514 127358
rect 115542 124978 115570 127414
rect 115710 126658 115738 130060
rect 115710 126625 115738 126630
rect 115934 128954 115962 128959
rect 115542 124950 115724 124978
rect 115934 124964 115962 128926
rect 116158 127498 116186 127503
rect 116158 124964 116186 127470
rect 116382 126546 116410 130060
rect 116886 128674 116914 128679
rect 116830 128170 116858 128175
rect 116382 126513 116410 126518
rect 116606 128114 116634 128119
rect 116382 126434 116410 126439
rect 116382 124964 116410 126406
rect 116606 124964 116634 128086
rect 116830 124964 116858 128142
rect 116886 124978 116914 128646
rect 117054 128618 117082 130060
rect 117726 128898 117754 130060
rect 117726 128865 117754 128870
rect 118398 128842 118426 130060
rect 119014 130046 119084 130074
rect 119518 130046 119756 130074
rect 118398 128809 118426 128814
rect 118622 129290 118650 129295
rect 117054 128585 117082 128590
rect 117502 126826 117530 126831
rect 117278 126434 117306 126439
rect 116886 124950 117068 124978
rect 117278 124964 117306 126406
rect 117502 124964 117530 126798
rect 118174 126658 118202 126663
rect 117726 126602 117754 126607
rect 117726 124964 117754 126574
rect 117950 126602 117978 126607
rect 117950 124964 117978 126574
rect 118174 124964 118202 126630
rect 118398 126546 118426 126551
rect 118398 124964 118426 126518
rect 118622 124964 118650 129262
rect 118846 128898 118874 128903
rect 118846 124964 118874 128870
rect 119014 126490 119042 130046
rect 119294 129178 119322 129183
rect 119014 126457 119042 126462
rect 119070 128842 119098 128847
rect 119070 124964 119098 128814
rect 119294 124964 119322 129150
rect 119518 124964 119546 130046
rect 120190 126938 120218 126943
rect 119742 126882 119770 126887
rect 119742 124964 119770 126854
rect 119966 126714 119994 126719
rect 119966 124964 119994 126686
rect 120190 124964 120218 126910
rect 120414 126882 120442 130060
rect 121086 129066 121114 130060
rect 121086 129033 121114 129038
rect 121310 129234 121338 129239
rect 120638 128898 120666 128903
rect 120414 126849 120442 126854
rect 120526 128562 120554 128567
rect 120526 124978 120554 128534
rect 120428 124950 120554 124978
rect 120638 124964 120666 128870
rect 121310 124964 121338 129206
rect 121758 126938 121786 130060
rect 121758 126905 121786 126910
rect 121982 129122 122010 129127
rect 121982 124964 122010 129094
rect 122430 128562 122458 130060
rect 123102 129010 123130 130060
rect 123102 128977 123130 128982
rect 123774 128954 123802 130060
rect 123774 128921 123802 128926
rect 122430 128529 122458 128534
rect 124446 128114 124474 130060
rect 124446 128081 124474 128086
rect 124670 129346 124698 129351
rect 122654 126658 122682 126663
rect 122654 124964 122682 126630
rect 123326 126546 123354 126551
rect 123326 124964 123354 126518
rect 123998 126490 124026 126495
rect 123998 124964 124026 126462
rect 124670 124964 124698 129318
rect 125118 126434 125146 130060
rect 125790 126602 125818 130060
rect 126462 129290 126490 130060
rect 126462 129257 126490 129262
rect 126686 129290 126714 129295
rect 125790 126569 125818 126574
rect 126014 129066 126042 129071
rect 125118 126401 125146 126406
rect 125342 126434 125370 126439
rect 125342 124964 125370 126406
rect 126014 124964 126042 129038
rect 126686 124964 126714 129262
rect 127134 129178 127162 130060
rect 127134 129145 127162 129150
rect 127358 129010 127386 129015
rect 127358 124964 127386 128982
rect 127806 126714 127834 130060
rect 128478 128898 128506 130060
rect 129150 129234 129178 130060
rect 129150 129201 129178 129206
rect 129822 129122 129850 130060
rect 129822 129089 129850 129094
rect 128478 128865 128506 128870
rect 127806 126681 127834 126686
rect 130494 126658 130522 130060
rect 130494 126625 130522 126630
rect 131166 126602 131194 130060
rect 131166 126569 131194 126574
rect 131838 126490 131866 130060
rect 132510 129346 132538 130060
rect 132510 129313 132538 129318
rect 131838 126457 131866 126462
rect 132286 128954 132314 128959
rect 78750 106521 78778 106526
rect 81550 106666 81578 106671
rect 79646 106498 79674 106503
rect 79646 104972 79674 106470
rect 81550 104972 81578 106638
rect 87262 106554 87290 106559
rect 83454 106386 83482 106391
rect 83454 104972 83482 106358
rect 85358 106330 85386 106335
rect 85358 104972 85386 106302
rect 87262 104972 87290 106526
rect 91070 106442 91098 106447
rect 89166 106274 89194 106279
rect 89166 104972 89194 106246
rect 91070 104972 91098 106414
rect 19278 75362 19306 75367
rect 19278 75329 19306 75334
rect 19278 75138 19306 75143
rect 18620 75054 18914 75082
rect 18886 74746 18914 75054
rect 16142 73738 16170 73743
rect 14294 73682 14322 73687
rect 13286 73626 13314 73631
rect 10430 73570 10458 73575
rect 9478 73514 9506 73519
rect 7574 7154 7602 7159
rect 6678 2170 6706 2175
rect 5782 2114 5810 2119
rect 5782 240 5810 2086
rect 6678 240 6706 2142
rect 7574 240 7602 7126
rect 8638 2954 8666 2959
rect 8638 240 8666 2926
rect 5684 196 5810 240
rect 5684 -480 5796 196
rect 6636 -480 6748 240
rect 7574 196 7700 240
rect 7588 -480 7700 196
rect 8540 196 8666 240
rect 9478 240 9506 73486
rect 10430 240 10458 73542
rect 12446 3010 12474 3015
rect 11494 2226 11522 2231
rect 11494 240 11522 2198
rect 12446 240 12474 2982
rect 9478 196 9604 240
rect 10430 196 10556 240
rect 8540 -480 8652 196
rect 9492 -480 9604 196
rect 10444 -480 10556 196
rect 11396 196 11522 240
rect 12348 196 12474 240
rect 13286 240 13314 73598
rect 14294 240 14322 73654
rect 15302 3066 15330 3071
rect 15302 240 15330 3038
rect 13286 196 13412 240
rect 11396 -480 11508 196
rect 12348 -480 12460 196
rect 13300 -480 13412 196
rect 14252 -480 14364 240
rect 15204 196 15330 240
rect 16142 240 16170 73710
rect 18494 73122 18522 73127
rect 18158 3178 18186 3183
rect 17206 3122 17234 3127
rect 17206 240 17234 3094
rect 18158 240 18186 3150
rect 18494 2170 18522 73094
rect 18494 2137 18522 2142
rect 18886 2114 18914 74718
rect 19278 73122 19306 75110
rect 19278 73089 19306 73094
rect 19950 7154 19978 75068
rect 19950 7121 19978 7126
rect 20622 2954 20650 75068
rect 21294 73514 21322 75068
rect 21966 73570 21994 75068
rect 21966 73537 21994 73542
rect 21294 73481 21322 73486
rect 21854 73514 21882 73519
rect 20622 2921 20650 2926
rect 20958 2394 20986 2399
rect 20062 2170 20090 2175
rect 18886 2081 18914 2086
rect 19110 2114 19138 2119
rect 19110 240 19138 2086
rect 20062 240 20090 2142
rect 20958 240 20986 2366
rect 21854 240 21882 73486
rect 22638 2226 22666 75068
rect 23310 3010 23338 75068
rect 23982 73626 24010 75068
rect 24654 73682 24682 75068
rect 24654 73649 24682 73654
rect 23982 73593 24010 73598
rect 24766 73626 24794 73631
rect 23310 2977 23338 2982
rect 23926 73570 23954 73575
rect 22638 2193 22666 2198
rect 22918 2170 22946 2175
rect 22918 240 22946 2142
rect 23926 2170 23954 73542
rect 24038 73178 24066 73183
rect 24038 2282 24066 73150
rect 24038 2249 24066 2254
rect 23926 2137 23954 2142
rect 23870 2058 23898 2063
rect 23870 240 23898 2030
rect 24766 2058 24794 73598
rect 24878 73122 24906 73127
rect 24878 2394 24906 73094
rect 25326 3066 25354 75068
rect 25998 73738 26026 75068
rect 25998 73705 26026 73710
rect 26446 73794 26474 73799
rect 25326 3033 25354 3038
rect 24878 2361 24906 2366
rect 24766 2025 24794 2030
rect 24822 2226 24850 2231
rect 24822 240 24850 2198
rect 26446 2226 26474 73766
rect 26670 3122 26698 75068
rect 27342 3178 27370 75068
rect 27342 3145 27370 3150
rect 26670 3089 26698 3094
rect 27678 2282 27706 2287
rect 26446 2193 26474 2198
rect 26726 2226 26754 2231
rect 25774 2170 25802 2175
rect 25774 240 25802 2142
rect 26726 240 26754 2198
rect 27678 240 27706 2254
rect 28014 2114 28042 75068
rect 28014 2081 28042 2086
rect 28574 73682 28602 73687
rect 28574 240 28602 73654
rect 28686 73178 28714 75068
rect 28686 73145 28714 73150
rect 29358 73122 29386 75068
rect 29358 73089 29386 73094
rect 29470 73738 29498 73743
rect 29470 240 29498 73710
rect 30030 73514 30058 75068
rect 30702 73570 30730 75068
rect 31374 73626 31402 75068
rect 32046 73794 32074 75068
rect 32046 73761 32074 73766
rect 31374 73593 31402 73598
rect 30702 73537 30730 73542
rect 30030 73481 30058 73486
rect 30422 73514 30450 73519
rect 30422 240 30450 73486
rect 32438 2338 32466 2343
rect 31486 2114 31514 2119
rect 31486 240 31514 2086
rect 32438 240 32466 2310
rect 32718 2170 32746 75068
rect 33390 4214 33418 75068
rect 33334 4186 33418 4214
rect 33334 2226 33362 4186
rect 34062 2394 34090 75068
rect 34734 73682 34762 75068
rect 35406 73738 35434 75068
rect 35406 73705 35434 73710
rect 34734 73649 34762 73654
rect 36078 73514 36106 75068
rect 36078 73481 36106 73486
rect 34062 2361 34090 2366
rect 34846 73122 34874 73127
rect 33334 2193 33362 2198
rect 33390 2282 33418 2287
rect 32718 2137 32746 2142
rect 33390 240 33418 2254
rect 34342 2114 34370 2119
rect 34342 240 34370 2086
rect 34846 2114 34874 73094
rect 36246 2450 36274 2455
rect 34846 2081 34874 2086
rect 35238 2114 35266 2119
rect 35238 240 35266 2086
rect 36246 240 36274 2422
rect 36750 2170 36778 75068
rect 36750 2137 36778 2142
rect 37198 2506 37226 2511
rect 37198 240 37226 2478
rect 37422 2338 37450 75068
rect 37422 2305 37450 2310
rect 38094 2282 38122 75068
rect 38766 73122 38794 75068
rect 38766 73089 38794 73094
rect 38990 73514 39018 73519
rect 38094 2249 38122 2254
rect 38150 2338 38178 2343
rect 38150 240 38178 2310
rect 16142 196 16268 240
rect 15204 -480 15316 196
rect 16156 -480 16268 196
rect 17108 196 17234 240
rect 18060 196 18186 240
rect 19012 196 19138 240
rect 19964 196 20090 240
rect 17108 -480 17220 196
rect 18060 -480 18172 196
rect 19012 -480 19124 196
rect 19964 -480 20076 196
rect 20916 -480 21028 240
rect 21854 196 21980 240
rect 21868 -480 21980 196
rect 22820 196 22946 240
rect 23772 196 23898 240
rect 24724 196 24850 240
rect 25676 196 25802 240
rect 26628 196 26754 240
rect 27580 196 27706 240
rect 22820 -480 22932 196
rect 23772 -480 23884 196
rect 24724 -480 24836 196
rect 25676 -480 25788 196
rect 26628 -480 26740 196
rect 27580 -480 27692 196
rect 28532 -480 28644 240
rect 29470 196 29596 240
rect 30422 196 30548 240
rect 29484 -480 29596 196
rect 30436 -480 30548 196
rect 31388 196 31514 240
rect 32340 196 32466 240
rect 33292 196 33418 240
rect 34244 196 34370 240
rect 31388 -480 31500 196
rect 32340 -480 32452 196
rect 33292 -480 33404 196
rect 34244 -480 34356 196
rect 35196 -480 35308 240
rect 36148 196 36274 240
rect 37100 196 37226 240
rect 38052 196 38178 240
rect 38990 240 39018 73486
rect 39438 2114 39466 75068
rect 40110 2450 40138 75068
rect 40782 2506 40810 75068
rect 40782 2473 40810 2478
rect 40110 2417 40138 2422
rect 41454 2338 41482 75068
rect 42126 73514 42154 75068
rect 42126 73481 42154 73486
rect 41454 2305 41482 2310
rect 41846 73178 41874 73183
rect 41006 2170 41034 2175
rect 39438 2081 39466 2086
rect 40054 2114 40082 2119
rect 40054 240 40082 2086
rect 41006 240 41034 2142
rect 38990 196 39116 240
rect 36148 -480 36260 196
rect 37100 -480 37212 196
rect 38052 -480 38164 196
rect 39004 -480 39116 196
rect 39956 196 40082 240
rect 40908 196 41034 240
rect 41846 240 41874 73150
rect 42798 2114 42826 75068
rect 43470 2170 43498 75068
rect 44142 73178 44170 75068
rect 44142 73145 44170 73150
rect 43470 2137 43498 2142
rect 43750 73122 43778 73127
rect 42798 2081 42826 2086
rect 42910 2114 42938 2119
rect 42910 240 42938 2086
rect 41846 196 41972 240
rect 39956 -480 40068 196
rect 40908 -480 41020 196
rect 41860 -480 41972 196
rect 42812 196 42938 240
rect 43750 240 43778 73094
rect 44814 4214 44842 75068
rect 45486 73122 45514 75068
rect 45486 73089 45514 73094
rect 44758 4186 44842 4214
rect 44758 2114 44786 4186
rect 44758 2081 44786 2086
rect 44814 2450 44842 2455
rect 44814 240 44842 2422
rect 46158 2450 46186 75068
rect 46158 2417 46186 2422
rect 45766 2170 45794 2175
rect 45766 240 45794 2142
rect 46830 2170 46858 75068
rect 46830 2137 46858 2142
rect 46718 2114 46746 2119
rect 46718 240 46746 2086
rect 47502 2114 47530 75068
rect 47502 2081 47530 2086
rect 47670 2114 47698 2119
rect 47670 240 47698 2086
rect 48174 2114 48202 75068
rect 48734 75054 48860 75082
rect 48734 73122 48762 75054
rect 49518 74774 49546 75068
rect 48174 2081 48202 2086
rect 48510 73094 48762 73122
rect 49462 74746 49546 74774
rect 43750 196 43876 240
rect 42812 -480 42924 196
rect 43764 -480 43876 196
rect 44716 196 44842 240
rect 45668 196 45794 240
rect 46620 196 46746 240
rect 47572 196 47698 240
rect 48510 240 48538 73094
rect 49462 240 49490 74746
rect 50190 2114 50218 75068
rect 50876 75054 51226 75082
rect 51198 73122 51226 75054
rect 51534 73122 51562 75068
rect 52206 73178 52234 75068
rect 52206 73145 52234 73150
rect 51198 73094 51282 73122
rect 51254 68894 51282 73094
rect 51534 73089 51562 73094
rect 52318 73122 52346 73127
rect 51254 68866 51394 68894
rect 50190 2086 50442 2114
rect 50414 240 50442 2086
rect 51366 240 51394 68866
rect 52318 240 52346 73094
rect 52878 73122 52906 75068
rect 52878 73089 52906 73094
rect 53270 73178 53298 73183
rect 53270 240 53298 73150
rect 53550 73178 53578 75068
rect 54222 73290 54250 75068
rect 54222 73257 54250 73262
rect 54894 73234 54922 75068
rect 54894 73201 54922 73206
rect 53550 73145 53578 73150
rect 55174 73178 55202 73183
rect 54166 73122 54194 73127
rect 54166 10094 54194 73094
rect 54166 10066 54250 10094
rect 54222 240 54250 10066
rect 55174 240 55202 73150
rect 55566 2506 55594 75068
rect 55566 2473 55594 2478
rect 56126 73290 56154 73295
rect 56126 240 56154 73262
rect 56238 2226 56266 75068
rect 56910 73570 56938 75068
rect 56910 73537 56938 73542
rect 56238 2193 56266 2198
rect 57134 73234 57162 73239
rect 57134 240 57162 73206
rect 57582 2114 57610 75068
rect 57582 2081 57610 2086
rect 58030 2506 58058 2511
rect 58030 240 58058 2478
rect 58254 2058 58282 75068
rect 58926 73122 58954 75068
rect 58926 73089 58954 73094
rect 59598 2506 59626 75068
rect 59598 2473 59626 2478
rect 59934 73570 59962 73575
rect 58254 2025 58282 2030
rect 58982 2226 59010 2231
rect 58982 240 59010 2198
rect 59934 240 59962 73542
rect 60270 2226 60298 75068
rect 60942 2282 60970 75068
rect 60942 2249 60970 2254
rect 60270 2193 60298 2198
rect 61614 2170 61642 75068
rect 62286 73626 62314 75068
rect 62286 73593 62314 73598
rect 62958 73514 62986 75068
rect 62958 73481 62986 73486
rect 61614 2137 61642 2142
rect 62790 73122 62818 73127
rect 60886 2114 60914 2119
rect 60886 240 60914 2086
rect 61838 2058 61866 2063
rect 61838 240 61866 2030
rect 62790 240 62818 73094
rect 63630 2058 63658 75068
rect 64302 73122 64330 75068
rect 64974 73234 65002 75068
rect 64974 73201 65002 73206
rect 65198 73626 65226 73631
rect 64302 73089 64330 73094
rect 65086 73122 65114 73127
rect 63630 2025 63658 2030
rect 63742 2506 63770 2511
rect 63742 240 63770 2478
rect 65086 2450 65114 73094
rect 65086 2417 65114 2422
rect 64694 2226 64722 2231
rect 64694 240 64722 2198
rect 65198 2114 65226 73598
rect 65646 73122 65674 75068
rect 66318 73178 66346 75068
rect 66990 73626 67018 75068
rect 66990 73593 67018 73598
rect 66318 73145 66346 73150
rect 65646 73089 65674 73094
rect 66766 73122 66794 73127
rect 65198 2081 65226 2086
rect 65646 2282 65674 2287
rect 65646 240 65674 2254
rect 66598 2170 66626 2175
rect 66598 240 66626 2142
rect 66766 2170 66794 73094
rect 67662 2282 67690 75068
rect 67662 2249 67690 2254
rect 67774 73514 67802 73519
rect 66766 2137 66794 2142
rect 67550 2114 67578 2119
rect 67550 240 67578 2086
rect 67774 2114 67802 73486
rect 68334 73514 68362 75068
rect 68334 73481 68362 73486
rect 68446 73178 68474 73183
rect 68446 2338 68474 73150
rect 69006 73122 69034 75068
rect 69006 73089 69034 73094
rect 69286 73234 69314 73239
rect 68446 2305 68474 2310
rect 67774 2081 67802 2086
rect 68502 2114 68530 2119
rect 68502 240 68530 2086
rect 69286 2058 69314 73206
rect 69678 3234 69706 75068
rect 69678 3201 69706 3206
rect 70350 3178 70378 75068
rect 70350 3145 70378 3150
rect 70966 73626 70994 73631
rect 70406 2450 70434 2455
rect 69286 2025 69314 2030
rect 69454 2114 69482 2119
rect 69454 240 69482 2086
rect 70406 240 70434 2422
rect 70966 2114 70994 73598
rect 71022 73178 71050 75068
rect 71022 73145 71050 73150
rect 71694 3122 71722 75068
rect 71694 3089 71722 3094
rect 72366 3066 72394 75068
rect 72366 3033 72394 3038
rect 72646 73514 72674 73519
rect 72646 2450 72674 73486
rect 72646 2417 72674 2422
rect 72758 73122 72786 73127
rect 72758 2226 72786 73094
rect 73038 73122 73066 75068
rect 73038 73089 73066 73094
rect 73486 73178 73514 73183
rect 72758 2193 72786 2198
rect 73262 2338 73290 2343
rect 70966 2081 70994 2086
rect 72310 2170 72338 2175
rect 71414 2058 71442 2063
rect 71414 240 71442 2030
rect 72310 240 72338 2142
rect 73262 240 73290 2310
rect 73486 2338 73514 73150
rect 73710 3010 73738 75068
rect 74382 73570 74410 75068
rect 74382 73537 74410 73542
rect 73710 2977 73738 2982
rect 73486 2305 73514 2310
rect 74214 2114 74242 2119
rect 74214 240 74242 2086
rect 75054 2114 75082 75068
rect 75166 73122 75194 73127
rect 75166 10094 75194 73094
rect 75166 10066 75250 10094
rect 75054 2081 75082 2086
rect 75166 2282 75194 2287
rect 75166 240 75194 2254
rect 75222 2170 75250 10066
rect 75726 3346 75754 75068
rect 75726 3313 75754 3318
rect 76398 2954 76426 75068
rect 77070 73626 77098 75068
rect 77070 73593 77098 73598
rect 77742 3290 77770 75068
rect 77742 3257 77770 3262
rect 76398 2921 76426 2926
rect 78022 3234 78050 3239
rect 75222 2137 75250 2142
rect 76118 2450 76146 2455
rect 76118 240 76146 2422
rect 77070 2226 77098 2231
rect 77070 240 77098 2198
rect 78022 240 78050 3206
rect 78414 2226 78442 75068
rect 79086 73738 79114 75068
rect 79086 73705 79114 73710
rect 79758 73122 79786 75068
rect 79758 73089 79786 73094
rect 80206 73122 80234 73127
rect 80206 3234 80234 73094
rect 80206 3201 80234 3206
rect 78414 2193 78442 2198
rect 78974 3178 79002 3183
rect 78974 240 79002 3150
rect 80430 3178 80458 75068
rect 81102 73514 81130 75068
rect 81102 73481 81130 73486
rect 80430 3145 80458 3150
rect 80878 3122 80906 3127
rect 79926 2338 79954 2343
rect 79926 240 79954 2310
rect 80878 240 80906 3094
rect 81774 3122 81802 75068
rect 82446 73850 82474 75068
rect 82446 73817 82474 73822
rect 81774 3089 81802 3094
rect 81830 3066 81858 3071
rect 81830 240 81858 3038
rect 82782 2170 82810 2175
rect 82782 240 82810 2142
rect 83118 2170 83146 75068
rect 83790 3066 83818 75068
rect 84462 73906 84490 75068
rect 84462 73873 84490 73878
rect 83790 3033 83818 3038
rect 84686 73570 84714 73575
rect 83118 2137 83146 2142
rect 83734 3010 83762 3015
rect 83734 240 83762 2982
rect 84686 240 84714 73542
rect 85134 73570 85162 75068
rect 85134 73537 85162 73542
rect 85806 3010 85834 75068
rect 85806 2977 85834 2982
rect 85694 2114 85722 2119
rect 85694 240 85722 2086
rect 86478 2114 86506 75068
rect 87150 73682 87178 75068
rect 87150 73649 87178 73654
rect 87766 73626 87794 73631
rect 86478 2081 86506 2086
rect 86590 3346 86618 3351
rect 86590 240 86618 3318
rect 87542 2954 87570 2959
rect 87542 240 87570 2926
rect 87766 2058 87794 73598
rect 87822 2954 87850 75068
rect 88494 73794 88522 75068
rect 88494 73761 88522 73766
rect 87822 2921 87850 2926
rect 88606 73738 88634 73743
rect 88606 2562 88634 73710
rect 89166 73626 89194 75068
rect 90286 73906 90314 73911
rect 89166 73593 89194 73598
rect 89502 73850 89530 73855
rect 88606 2529 88634 2534
rect 89446 3290 89474 3295
rect 87766 2025 87794 2030
rect 88494 2058 88522 2063
rect 88494 240 88522 2030
rect 89446 240 89474 3262
rect 89502 2338 89530 73822
rect 89502 2305 89530 2310
rect 90286 2282 90314 73878
rect 96166 73794 96194 73799
rect 93646 73514 93674 73519
rect 92302 3234 92330 3239
rect 90286 2249 90314 2254
rect 91350 2562 91378 2567
rect 90398 2226 90426 2231
rect 90398 240 90426 2198
rect 91350 240 91378 2534
rect 92302 240 92330 3206
rect 93254 3178 93282 3183
rect 93254 240 93282 3150
rect 93646 2170 93674 73486
rect 96166 10094 96194 73766
rect 97846 73682 97874 73687
rect 96278 73570 96306 73575
rect 96166 10066 96250 10094
rect 95158 3122 95186 3127
rect 93646 2137 93674 2142
rect 94206 2170 94234 2175
rect 94206 240 94234 2142
rect 95158 240 95186 3094
rect 96110 2338 96138 2343
rect 96110 240 96138 2310
rect 96222 2338 96250 10066
rect 96278 2394 96306 73542
rect 96278 2361 96306 2366
rect 96222 2305 96250 2310
rect 97230 2338 97258 2343
rect 97230 2226 97258 2310
rect 97846 2338 97874 73654
rect 99526 73626 99554 73631
rect 97846 2305 97874 2310
rect 98014 3066 98042 3071
rect 97230 2193 97258 2198
rect 97062 2170 97090 2175
rect 97062 240 97090 2142
rect 98014 240 98042 3038
rect 98966 2282 98994 2287
rect 98966 240 98994 2254
rect 99526 2170 99554 73598
rect 100870 3010 100898 3015
rect 99526 2137 99554 2142
rect 99974 2394 100002 2399
rect 99974 240 100002 2366
rect 100870 240 100898 2982
rect 103726 2954 103754 2959
rect 102774 2338 102802 2343
rect 101822 2114 101850 2119
rect 101822 240 101850 2086
rect 102774 240 102802 2310
rect 103726 240 103754 2926
rect 104678 2226 104706 2231
rect 104678 240 104706 2198
rect 105630 2170 105658 2175
rect 105630 240 105658 2142
rect 129542 2114 129570 2119
rect 129542 240 129570 2086
rect 132286 240 132314 128926
rect 133182 126434 133210 130060
rect 133854 129066 133882 130060
rect 134526 129290 134554 130060
rect 134526 129257 134554 129262
rect 133854 129033 133882 129038
rect 135198 129010 135226 130060
rect 135198 128977 135226 128982
rect 137998 129010 138026 129015
rect 133182 126401 133210 126406
rect 135198 2170 135226 2175
rect 135198 240 135226 2142
rect 137998 240 138026 128982
rect 142590 2114 142618 130060
rect 143262 128954 143290 130060
rect 143262 128921 143290 128926
rect 142590 2081 142618 2086
rect 143822 2506 143850 2511
rect 140966 2058 140994 2063
rect 140966 240 140994 2030
rect 143822 240 143850 2478
rect 143934 2170 143962 130060
rect 144606 129010 144634 130060
rect 144606 128977 144634 128982
rect 143934 2137 143962 2142
rect 145278 2058 145306 130060
rect 145950 2506 145978 130060
rect 145950 2473 145978 2478
rect 146566 130046 146636 130074
rect 145278 2025 145306 2030
rect 146566 240 146594 130046
rect 147294 2114 147322 130060
rect 147966 2450 147994 130060
rect 148638 129010 148666 130060
rect 148638 128977 148666 128982
rect 149310 2954 149338 130060
rect 149982 128954 150010 130060
rect 149982 128921 150010 128926
rect 149310 2921 149338 2926
rect 147966 2417 147994 2422
rect 150654 2282 150682 130060
rect 150654 2249 150682 2254
rect 151326 2226 151354 130060
rect 151326 2193 151354 2198
rect 151998 2170 152026 130060
rect 151998 2137 152026 2142
rect 152278 2450 152306 2455
rect 147294 2081 147322 2086
rect 149422 2114 149450 2119
rect 149422 240 149450 2086
rect 152278 240 152306 2422
rect 152670 2114 152698 130060
rect 172102 129122 172130 129127
rect 170982 129066 171010 129071
rect 152670 2081 152698 2086
rect 155134 129010 155162 129015
rect 155134 240 155162 128982
rect 169862 129010 169890 129015
rect 159166 128954 159194 128959
rect 157990 2954 158018 2959
rect 157990 240 158018 2926
rect 159166 2058 159194 128926
rect 163142 128954 163170 128959
rect 163142 124964 163170 128926
rect 168742 126546 168770 126551
rect 167622 126490 167650 126495
rect 166502 126434 166530 126439
rect 166502 124964 166530 126406
rect 167622 124964 167650 126462
rect 168742 124964 168770 126518
rect 169862 124964 169890 128982
rect 170982 124964 171010 129038
rect 172102 124964 172130 129094
rect 173502 128954 173530 130060
rect 173502 128921 173530 128926
rect 174342 128954 174370 128959
rect 173222 126602 173250 126607
rect 173222 124964 173250 126574
rect 174342 124964 174370 128926
rect 175462 128114 175490 128119
rect 175462 124964 175490 128086
rect 175518 126434 175546 130060
rect 176190 126490 176218 130060
rect 176190 126457 176218 126462
rect 176582 126826 176610 126831
rect 175518 126401 175546 126406
rect 176582 124964 176610 126798
rect 176862 126546 176890 130060
rect 177534 129010 177562 130060
rect 178206 129066 178234 130060
rect 178878 129122 178906 130060
rect 178878 129089 178906 129094
rect 178206 129033 178234 129038
rect 178822 129066 178850 129071
rect 177534 128977 177562 128982
rect 176862 126513 176890 126518
rect 177702 128562 177730 128567
rect 177702 124964 177730 128534
rect 178822 124964 178850 129038
rect 179550 126602 179578 130060
rect 179550 126569 179578 126574
rect 179942 129122 179970 129127
rect 179942 124964 179970 129094
rect 180222 128954 180250 130060
rect 180222 128921 180250 128926
rect 180894 128114 180922 130060
rect 180894 128081 180922 128086
rect 181062 128898 181090 128903
rect 181062 124964 181090 128870
rect 181566 126826 181594 130060
rect 181566 126793 181594 126798
rect 182182 128954 182210 128959
rect 182182 124964 182210 128926
rect 182238 128562 182266 130060
rect 182910 129066 182938 130060
rect 183582 129122 183610 130060
rect 183582 129089 183610 129094
rect 182910 129033 182938 129038
rect 184254 128898 184282 130060
rect 184926 128954 184954 130060
rect 184926 128921 184954 128926
rect 184254 128865 184282 128870
rect 184422 128898 184450 128903
rect 182238 128529 182266 128534
rect 183302 128842 183330 128847
rect 183302 124964 183330 128814
rect 184422 124964 184450 128870
rect 185598 128842 185626 130060
rect 186270 128898 186298 130060
rect 186270 128865 186298 128870
rect 185598 128809 185626 128814
rect 185542 128562 185570 128567
rect 185542 124964 185570 128534
rect 186942 128562 186970 130060
rect 186942 128529 186970 128534
rect 186662 126882 186690 126887
rect 186662 124964 186690 126854
rect 187614 126882 187642 130060
rect 188286 127694 188314 130060
rect 187614 126849 187642 126854
rect 188118 127666 188314 127694
rect 188902 130046 188972 130074
rect 189644 130046 189826 130074
rect 188118 124978 188146 127666
rect 187796 124950 188146 124978
rect 188902 124964 188930 130046
rect 189798 128898 189826 130046
rect 190302 128898 190330 130060
rect 189798 128870 189882 128898
rect 189854 124978 189882 128870
rect 190302 128865 190330 128870
rect 190974 128842 191002 130060
rect 190974 128809 191002 128814
rect 191142 128898 191170 128903
rect 189854 124950 190036 124978
rect 191142 124964 191170 128870
rect 191646 126826 191674 130060
rect 191646 126793 191674 126798
rect 192262 128842 192290 128847
rect 192262 124964 192290 128814
rect 192318 126434 192346 130060
rect 192318 126401 192346 126406
rect 192990 126266 193018 130060
rect 192990 126233 193018 126238
rect 193382 126826 193410 126831
rect 193382 124964 193410 126798
rect 193662 126210 193690 130060
rect 193662 126177 193690 126182
rect 194334 126154 194362 130060
rect 195006 126770 195034 130060
rect 195678 129066 195706 130060
rect 195678 129033 195706 129038
rect 196350 129010 196378 130060
rect 196350 128977 196378 128982
rect 197022 128954 197050 130060
rect 197022 128921 197050 128926
rect 197694 128170 197722 130060
rect 197694 128137 197722 128142
rect 198366 128114 198394 130060
rect 198366 128081 198394 128086
rect 195006 126737 195034 126742
rect 198982 126770 199010 126775
rect 194334 126121 194362 126126
rect 194502 126434 194530 126439
rect 194502 124964 194530 126406
rect 195622 126266 195650 126271
rect 195622 124964 195650 126238
rect 196742 126210 196770 126215
rect 196742 124964 196770 126182
rect 197862 126154 197890 126159
rect 197862 124964 197890 126126
rect 198982 124964 199010 126742
rect 199038 126714 199066 130060
rect 199710 127330 199738 130060
rect 199710 127297 199738 127302
rect 200102 129066 200130 129071
rect 199038 126681 199066 126686
rect 200102 124964 200130 129038
rect 200382 126658 200410 130060
rect 200382 126625 200410 126630
rect 201054 126602 201082 130060
rect 201054 126569 201082 126574
rect 201222 129010 201250 129015
rect 201222 124964 201250 128982
rect 201726 127274 201754 130060
rect 201726 127241 201754 127246
rect 202342 128954 202370 128959
rect 202342 124964 202370 128926
rect 202398 126546 202426 130060
rect 203070 127554 203098 130060
rect 203742 129122 203770 130060
rect 203742 129089 203770 129094
rect 204414 128954 204442 130060
rect 204414 128921 204442 128926
rect 203070 127521 203098 127526
rect 203462 128170 203490 128175
rect 202398 126513 202426 126518
rect 203462 124964 203490 128142
rect 204582 128114 204610 128119
rect 204582 124964 204610 128086
rect 205086 126490 205114 130060
rect 205086 126457 205114 126462
rect 205702 126714 205730 126719
rect 205702 124964 205730 126686
rect 205758 126434 205786 130060
rect 205758 126401 205786 126406
rect 206430 126378 206458 130060
rect 206430 126345 206458 126350
rect 206822 127330 206850 127335
rect 206822 124964 206850 127302
rect 207102 126826 207130 130060
rect 207774 127498 207802 130060
rect 207774 127465 207802 127470
rect 208446 127442 208474 130060
rect 208446 127409 208474 127414
rect 209118 127386 209146 130060
rect 209118 127353 209146 127358
rect 209790 127330 209818 130060
rect 210462 129066 210490 130060
rect 210462 129033 210490 129038
rect 209790 127297 209818 127302
rect 207102 126793 207130 126798
rect 210182 127274 210210 127279
rect 207942 126658 207970 126663
rect 207942 124964 207970 126630
rect 209062 126602 209090 126607
rect 209062 124964 209090 126574
rect 210182 124964 210210 127246
rect 211134 127274 211162 130060
rect 211806 129010 211834 130060
rect 211806 128977 211834 128982
rect 212478 128114 212506 130060
rect 212478 128081 212506 128086
rect 211134 127241 211162 127246
rect 212422 127554 212450 127559
rect 211302 126546 211330 126551
rect 211302 124964 211330 126518
rect 212422 124964 212450 127526
rect 213150 126770 213178 130060
rect 213150 126737 213178 126742
rect 213542 129122 213570 129127
rect 213542 124964 213570 129094
rect 213822 126714 213850 130060
rect 213822 126681 213850 126686
rect 214494 126658 214522 130060
rect 214494 126625 214522 126630
rect 214662 128954 214690 128959
rect 214662 124964 214690 128926
rect 215166 126602 215194 130060
rect 215166 126569 215194 126574
rect 215838 126546 215866 130060
rect 215838 126513 215866 126518
rect 215782 126490 215810 126495
rect 215782 124964 215810 126462
rect 216510 126490 216538 130060
rect 216510 126457 216538 126462
rect 216902 126434 216930 126439
rect 216902 124964 216930 126406
rect 217182 126434 217210 130060
rect 217854 128954 217882 130060
rect 222558 129122 222586 130060
rect 223230 129234 223258 130060
rect 223230 129201 223258 129206
rect 222558 129089 222586 129094
rect 217854 128921 217882 128926
rect 223902 128562 223930 130060
rect 224574 129178 224602 130060
rect 224574 129145 224602 129150
rect 223902 128529 223930 128534
rect 224742 129066 224770 129071
rect 220262 127498 220290 127503
rect 217182 126401 217210 126406
rect 219142 126826 219170 126831
rect 218022 126378 218050 126383
rect 218022 124964 218050 126350
rect 219142 124964 219170 126798
rect 220262 124964 220290 127470
rect 221382 127442 221410 127447
rect 221382 124964 221410 127414
rect 222502 127386 222530 127391
rect 222502 124964 222530 127358
rect 223622 127330 223650 127335
rect 223622 124964 223650 127302
rect 224742 124964 224770 129038
rect 225246 127554 225274 130060
rect 225246 127521 225274 127526
rect 225862 127274 225890 127279
rect 225862 124964 225890 127246
rect 225918 126826 225946 130060
rect 226590 127498 226618 130060
rect 226590 127465 226618 127470
rect 226982 129010 227010 129015
rect 225918 126793 225946 126798
rect 226982 124964 227010 128982
rect 227262 127442 227290 130060
rect 227262 127409 227290 127414
rect 227934 127386 227962 130060
rect 228494 128562 228522 128567
rect 227934 127353 227962 127358
rect 228102 128114 228130 128119
rect 228102 124964 228130 128086
rect 228494 126378 228522 128534
rect 228606 127330 228634 130060
rect 228606 127297 228634 127302
rect 229278 127274 229306 130060
rect 229950 128338 229978 130060
rect 229950 128305 229978 128310
rect 230622 128282 230650 130060
rect 230622 128249 230650 128254
rect 230958 129234 230986 129239
rect 229278 127241 229306 127246
rect 228494 126345 228522 126350
rect 229222 126770 229250 126775
rect 229222 124964 229250 126742
rect 230342 126714 230370 126719
rect 230342 124964 230370 126686
rect 230958 126266 230986 129206
rect 231294 128226 231322 130060
rect 231294 128193 231322 128198
rect 231798 129122 231826 129127
rect 230958 126233 230986 126238
rect 231462 126658 231490 126663
rect 231462 124964 231490 126630
rect 231798 126658 231826 129094
rect 231966 128170 231994 130060
rect 231966 128137 231994 128142
rect 232246 129178 232274 129183
rect 231798 126625 231826 126630
rect 232246 126322 232274 129150
rect 232638 129010 232666 130060
rect 233310 129290 233338 130060
rect 233310 129257 233338 129262
rect 233982 129234 234010 130060
rect 233982 129201 234010 129206
rect 234654 129122 234682 130060
rect 234654 129089 234682 129094
rect 232638 128977 232666 128982
rect 233814 128954 233842 128959
rect 232246 126289 232274 126294
rect 232582 126602 232610 126607
rect 232582 124964 232610 126574
rect 233702 126546 233730 126551
rect 233702 124964 233730 126518
rect 233814 126210 233842 128926
rect 235326 128114 235354 130060
rect 235998 129066 236026 130060
rect 236670 129346 236698 130060
rect 236670 129313 236698 129318
rect 235998 129033 236026 129038
rect 237342 128954 237370 130060
rect 237342 128921 237370 128926
rect 235326 128081 235354 128086
rect 238014 126770 238042 130060
rect 238014 126737 238042 126742
rect 238686 126714 238714 130060
rect 238686 126681 238714 126686
rect 238182 126658 238210 126663
rect 233814 126177 233842 126182
rect 234822 126490 234850 126495
rect 234822 124964 234850 126462
rect 235942 126434 235970 126439
rect 235942 124964 235970 126406
rect 237062 126210 237090 126215
rect 237062 124964 237090 126182
rect 238182 124964 238210 126630
rect 239358 126658 239386 130060
rect 239414 129010 239442 129015
rect 239414 127610 239442 128982
rect 240030 129010 240058 130060
rect 240030 128977 240058 128982
rect 239414 127577 239442 127582
rect 239358 126625 239386 126630
rect 240702 126602 240730 130060
rect 241374 129178 241402 130060
rect 241374 129145 241402 129150
rect 240702 126569 240730 126574
rect 242046 126546 242074 130060
rect 242046 126513 242074 126518
rect 242606 130046 242732 130074
rect 242606 126490 242634 130046
rect 242718 129290 242746 129295
rect 242718 127666 242746 129262
rect 242718 127633 242746 127638
rect 242606 126457 242634 126462
rect 242662 127554 242690 127559
rect 240422 126378 240450 126383
rect 239302 126266 239330 126271
rect 239302 124964 239330 126238
rect 240422 124964 240450 126350
rect 241542 126322 241570 126327
rect 241542 124964 241570 126294
rect 242662 124964 242690 127526
rect 243390 126434 243418 130060
rect 245014 129346 245042 129351
rect 243558 129234 243586 129239
rect 243558 127554 243586 129206
rect 243558 127521 243586 127526
rect 244902 127498 244930 127503
rect 243390 126401 243418 126406
rect 243782 126826 243810 126831
rect 243782 124964 243810 126798
rect 244902 124964 244930 127470
rect 245014 127498 245042 129318
rect 251566 129178 251594 129183
rect 245014 127465 245042 127470
rect 250502 128506 250530 128511
rect 246022 127442 246050 127447
rect 246022 124964 246050 127414
rect 247142 127386 247170 127391
rect 247142 124964 247170 127358
rect 248262 127330 248290 127335
rect 248262 124964 248290 127302
rect 249382 127274 249410 127279
rect 249382 124964 249410 127246
rect 250502 124964 250530 128478
rect 251566 128282 251594 129150
rect 258342 129122 258370 129127
rect 251566 128249 251594 128254
rect 251622 128450 251650 128455
rect 251622 124964 251650 128422
rect 252742 128170 252770 128175
rect 252742 124964 252770 128142
rect 253862 128058 253890 128063
rect 253862 124964 253890 128030
rect 256102 127666 256130 127671
rect 254982 127610 255010 127615
rect 254982 124964 255010 127582
rect 256102 124964 256130 127638
rect 257222 127554 257250 127559
rect 257222 124964 257250 127526
rect 258342 124964 258370 129094
rect 260582 129066 260610 129071
rect 259462 128114 259490 128119
rect 259462 124964 259490 128086
rect 260582 124964 260610 129038
rect 265398 129010 265426 129015
rect 262822 128954 262850 128959
rect 261702 127498 261730 127503
rect 261702 124964 261730 127470
rect 262822 124964 262850 128926
rect 263942 126770 263970 126775
rect 263942 124964 263970 126742
rect 265062 126714 265090 126719
rect 265062 124964 265090 126686
rect 265398 126210 265426 128982
rect 269542 128282 269570 128287
rect 265398 126177 265426 126182
rect 266182 126658 266210 126663
rect 266182 124964 266210 126630
rect 268422 126602 268450 126607
rect 267302 126210 267330 126215
rect 267302 124964 267330 126182
rect 268422 124964 268450 126574
rect 269542 124964 269570 128254
rect 270662 126546 270690 126551
rect 270662 124964 270690 126518
rect 271782 126490 271810 126495
rect 271782 124964 271810 126462
rect 272118 124810 272146 135254
rect 272902 126434 272930 126439
rect 272902 124964 272930 126406
rect 272118 124777 272146 124782
rect 269374 7154 269402 7159
rect 260806 6426 260834 6431
rect 249382 6370 249410 6375
rect 243670 6314 243698 6319
rect 163702 2282 163730 2287
rect 159166 2025 159194 2030
rect 160846 2058 160874 2063
rect 160846 240 160874 2030
rect 163702 240 163730 2254
rect 166558 2226 166586 2231
rect 166558 240 166586 2198
rect 169414 2170 169442 2175
rect 169414 240 169442 2142
rect 172270 2114 172298 2119
rect 172270 240 172298 2086
rect 243670 240 243698 6286
rect 246638 3794 246666 3799
rect 246638 240 246666 3766
rect 249382 240 249410 6342
rect 252350 4634 252378 4639
rect 252350 240 252378 4606
rect 255206 3850 255234 3855
rect 255206 240 255234 3822
rect 258062 2954 258090 2959
rect 258062 240 258090 2926
rect 260806 240 260834 6398
rect 266630 3066 266658 3071
rect 263718 3010 263746 3015
rect 263718 240 263746 2982
rect 266630 240 266658 3038
rect 269374 240 269402 7126
rect 272342 2114 272370 2119
rect 272342 240 272370 2086
rect 275198 240 275282 266
rect 48510 196 48636 240
rect 49462 196 49588 240
rect 50414 196 50540 240
rect 51366 196 51492 240
rect 52318 196 52444 240
rect 53270 196 53396 240
rect 54222 196 54348 240
rect 55174 196 55300 240
rect 56126 196 56252 240
rect 44716 -480 44828 196
rect 45668 -480 45780 196
rect 46620 -480 46732 196
rect 47572 -480 47684 196
rect 48524 -480 48636 196
rect 49476 -480 49588 196
rect 50428 -480 50540 196
rect 51380 -480 51492 196
rect 52332 -480 52444 196
rect 53284 -480 53396 196
rect 54236 -480 54348 196
rect 55188 -480 55300 196
rect 56140 -480 56252 196
rect 57092 -480 57204 240
rect 58030 196 58156 240
rect 58982 196 59108 240
rect 59934 196 60060 240
rect 60886 196 61012 240
rect 61838 196 61964 240
rect 62790 196 62916 240
rect 63742 196 63868 240
rect 64694 196 64820 240
rect 65646 196 65772 240
rect 66598 196 66724 240
rect 67550 196 67676 240
rect 68502 196 68628 240
rect 69454 196 69580 240
rect 70406 196 70532 240
rect 58044 -480 58156 196
rect 58996 -480 59108 196
rect 59948 -480 60060 196
rect 60900 -480 61012 196
rect 61852 -480 61964 196
rect 62804 -480 62916 196
rect 63756 -480 63868 196
rect 64708 -480 64820 196
rect 65660 -480 65772 196
rect 66612 -480 66724 196
rect 67564 -480 67676 196
rect 68516 -480 68628 196
rect 69468 -480 69580 196
rect 70420 -480 70532 196
rect 71372 -480 71484 240
rect 72310 196 72436 240
rect 73262 196 73388 240
rect 74214 196 74340 240
rect 75166 196 75292 240
rect 76118 196 76244 240
rect 77070 196 77196 240
rect 78022 196 78148 240
rect 78974 196 79100 240
rect 79926 196 80052 240
rect 80878 196 81004 240
rect 81830 196 81956 240
rect 82782 196 82908 240
rect 83734 196 83860 240
rect 84686 196 84812 240
rect 72324 -480 72436 196
rect 73276 -480 73388 196
rect 74228 -480 74340 196
rect 75180 -480 75292 196
rect 76132 -480 76244 196
rect 77084 -480 77196 196
rect 78036 -480 78148 196
rect 78988 -480 79100 196
rect 79940 -480 80052 196
rect 80892 -480 81004 196
rect 81844 -480 81956 196
rect 82796 -480 82908 196
rect 83748 -480 83860 196
rect 84700 -480 84812 196
rect 85652 -480 85764 240
rect 86590 196 86716 240
rect 87542 196 87668 240
rect 88494 196 88620 240
rect 89446 196 89572 240
rect 90398 196 90524 240
rect 91350 196 91476 240
rect 92302 196 92428 240
rect 93254 196 93380 240
rect 94206 196 94332 240
rect 95158 196 95284 240
rect 96110 196 96236 240
rect 97062 196 97188 240
rect 98014 196 98140 240
rect 98966 196 99092 240
rect 86604 -480 86716 196
rect 87556 -480 87668 196
rect 88508 -480 88620 196
rect 89460 -480 89572 196
rect 90412 -480 90524 196
rect 91364 -480 91476 196
rect 92316 -480 92428 196
rect 93268 -480 93380 196
rect 94220 -480 94332 196
rect 95172 -480 95284 196
rect 96124 -480 96236 196
rect 97076 -480 97188 196
rect 98028 -480 98140 196
rect 98980 -480 99092 196
rect 99932 -480 100044 240
rect 100870 196 100996 240
rect 101822 196 101948 240
rect 102774 196 102900 240
rect 103726 196 103852 240
rect 104678 196 104804 240
rect 105630 196 105756 240
rect 100884 -480 100996 196
rect 101836 -480 101948 196
rect 102788 -480 102900 196
rect 103740 -480 103852 196
rect 104692 -480 104804 196
rect 105644 -480 105756 196
rect 106596 -480 106708 240
rect 107548 -480 107660 240
rect 108500 -480 108612 240
rect 109452 -480 109564 240
rect 110404 -480 110516 240
rect 111356 -480 111468 240
rect 112308 -480 112420 240
rect 113260 -480 113372 240
rect 114212 -480 114324 240
rect 115164 -480 115276 240
rect 116116 -480 116228 240
rect 117068 -480 117180 240
rect 118020 -480 118132 240
rect 118972 -480 119084 240
rect 119924 -480 120036 240
rect 120876 -480 120988 240
rect 121828 -480 121940 240
rect 122780 -480 122892 240
rect 123732 -480 123844 240
rect 124684 -480 124796 240
rect 125636 -480 125748 240
rect 126588 -480 126700 240
rect 127540 -480 127652 240
rect 128492 -480 128604 240
rect 129444 196 129570 240
rect 129444 -480 129556 196
rect 130396 -480 130508 240
rect 131348 -480 131460 240
rect 132286 196 132412 240
rect 132300 -480 132412 196
rect 133252 -480 133364 240
rect 134204 -480 134316 240
rect 135156 -480 135268 240
rect 136108 -480 136220 240
rect 137060 -480 137172 240
rect 137998 196 138124 240
rect 138012 -480 138124 196
rect 138964 -480 139076 240
rect 139916 -480 140028 240
rect 140868 196 140994 240
rect 140868 -480 140980 196
rect 141820 -480 141932 240
rect 142772 -480 142884 240
rect 143724 196 143850 240
rect 143724 -480 143836 196
rect 144676 -480 144788 240
rect 145628 -480 145740 240
rect 146566 196 146692 240
rect 146580 -480 146692 196
rect 147532 -480 147644 240
rect 148484 -480 148596 240
rect 149422 196 149548 240
rect 149436 -480 149548 196
rect 150388 -480 150500 240
rect 151340 -480 151452 240
rect 152278 196 152404 240
rect 152292 -480 152404 196
rect 153244 -480 153356 240
rect 154196 -480 154308 240
rect 155134 196 155260 240
rect 155148 -480 155260 196
rect 156100 -480 156212 240
rect 157052 -480 157164 240
rect 157990 196 158116 240
rect 158004 -480 158116 196
rect 158956 -480 159068 240
rect 159908 -480 160020 240
rect 160846 196 160972 240
rect 160860 -480 160972 196
rect 161812 -480 161924 240
rect 162764 -480 162876 240
rect 163702 196 163828 240
rect 163716 -480 163828 196
rect 164668 -480 164780 240
rect 165620 -480 165732 240
rect 166558 196 166684 240
rect 166572 -480 166684 196
rect 167524 -480 167636 240
rect 168476 -480 168588 240
rect 169414 196 169540 240
rect 169428 -480 169540 196
rect 170380 -480 170492 240
rect 171332 -480 171444 240
rect 172270 196 172396 240
rect 172284 -480 172396 196
rect 173236 -480 173348 240
rect 174188 -480 174300 240
rect 175140 -480 175252 240
rect 176092 -480 176204 240
rect 177044 -480 177156 240
rect 177996 -480 178108 240
rect 178948 -480 179060 240
rect 179900 -480 180012 240
rect 180852 -480 180964 240
rect 181804 -480 181916 240
rect 182756 -480 182868 240
rect 183708 -480 183820 240
rect 184660 -480 184772 240
rect 185612 -480 185724 240
rect 186564 -480 186676 240
rect 187516 -480 187628 240
rect 188468 -480 188580 240
rect 189420 -480 189532 240
rect 190372 -480 190484 240
rect 191324 -480 191436 240
rect 192276 -480 192388 240
rect 193228 -480 193340 240
rect 194180 -480 194292 240
rect 195132 -480 195244 240
rect 196084 -480 196196 240
rect 197036 -480 197148 240
rect 197988 -480 198100 240
rect 198940 -480 199052 240
rect 199892 -480 200004 240
rect 200844 -480 200956 240
rect 201796 -480 201908 240
rect 202748 -480 202860 240
rect 203700 -480 203812 240
rect 204652 -480 204764 240
rect 205604 -480 205716 240
rect 206556 -480 206668 240
rect 207508 -480 207620 240
rect 208460 -480 208572 240
rect 209412 -480 209524 240
rect 210364 -480 210476 240
rect 211316 -480 211428 240
rect 212268 -480 212380 240
rect 213220 -480 213332 240
rect 214172 -480 214284 240
rect 215124 -480 215236 240
rect 216076 -480 216188 240
rect 217028 -480 217140 240
rect 217980 -480 218092 240
rect 218932 -480 219044 240
rect 219884 -480 219996 240
rect 220836 -480 220948 240
rect 221788 -480 221900 240
rect 222740 -480 222852 240
rect 223692 -480 223804 240
rect 224644 -480 224756 240
rect 225596 -480 225708 240
rect 226548 -480 226660 240
rect 227500 -480 227612 240
rect 228452 -480 228564 240
rect 229404 -480 229516 240
rect 230356 -480 230468 240
rect 231308 -480 231420 240
rect 232260 -480 232372 240
rect 233212 -480 233324 240
rect 234164 -480 234276 240
rect 235116 -480 235228 240
rect 236068 -480 236180 240
rect 237020 -480 237132 240
rect 237972 -480 238084 240
rect 238924 -480 239036 240
rect 239876 -480 239988 240
rect 240828 -480 240940 240
rect 241780 -480 241892 240
rect 242732 -480 242844 240
rect 243670 196 243796 240
rect 243684 -480 243796 196
rect 244636 -480 244748 240
rect 245588 -480 245700 240
rect 246540 196 246666 240
rect 246540 -480 246652 196
rect 247492 -480 247604 240
rect 248444 -480 248556 240
rect 249382 196 249508 240
rect 249396 -480 249508 196
rect 250348 -480 250460 240
rect 251300 -480 251412 240
rect 252252 196 252378 240
rect 252252 -480 252364 196
rect 253204 -480 253316 240
rect 254156 -480 254268 240
rect 255108 196 255234 240
rect 255108 -480 255220 196
rect 256060 -480 256172 240
rect 257012 -480 257124 240
rect 257964 196 258090 240
rect 257964 -480 258076 196
rect 258916 -480 259028 240
rect 259868 -480 259980 240
rect 260806 196 260932 240
rect 260820 -480 260932 196
rect 261772 -480 261884 240
rect 262724 -480 262836 240
rect 263676 -480 263788 240
rect 264628 -480 264740 240
rect 265580 -480 265692 240
rect 266532 196 266658 240
rect 266532 -480 266644 196
rect 267484 -480 267596 240
rect 268436 -480 268548 240
rect 269374 196 269500 240
rect 269388 -480 269500 196
rect 270340 -480 270452 240
rect 271292 -480 271404 240
rect 272244 196 272370 240
rect 272244 -480 272356 196
rect 273196 -480 273308 240
rect 274148 -480 274260 240
rect 275100 238 275282 240
rect 275100 196 275226 238
rect 275254 210 275282 238
rect 275422 210 275450 135646
rect 276430 134386 276458 134391
rect 276374 133938 276402 133943
rect 275590 133042 275618 133047
rect 275590 2954 275618 133014
rect 275646 132594 275674 132599
rect 275646 3850 275674 132566
rect 275646 3817 275674 3822
rect 276374 3010 276402 133910
rect 276430 3066 276458 134358
rect 277214 131698 277242 131703
rect 276430 3033 276458 3038
rect 276486 124810 276514 124815
rect 276374 2977 276402 2982
rect 275590 2921 275618 2926
rect 276486 2114 276514 124782
rect 277214 6370 277242 131670
rect 277214 6337 277242 6342
rect 276486 2081 276514 2086
rect 277606 2114 277634 137494
rect 277718 137074 277746 137079
rect 277718 2170 277746 137046
rect 277830 136626 277858 136631
rect 277830 2506 277858 136598
rect 277830 2473 277858 2478
rect 277942 136178 277970 136183
rect 277718 2137 277746 2142
rect 277606 2081 277634 2086
rect 277942 240 277970 136150
rect 278166 134834 278194 134839
rect 278054 132146 278082 132151
rect 278054 4634 278082 132118
rect 278054 4601 278082 4606
rect 278110 131250 278138 131255
rect 278110 3794 278138 131222
rect 278166 7154 278194 134806
rect 278166 7121 278194 7126
rect 278222 133490 278250 133495
rect 278222 6426 278250 133462
rect 278222 6393 278250 6398
rect 278278 130802 278306 130807
rect 278278 6314 278306 130774
rect 278278 6281 278306 6286
rect 278110 3761 278138 3766
rect 280798 2506 280826 2511
rect 280798 240 280826 2478
rect 283654 2170 283682 2175
rect 283654 240 283682 2142
rect 286510 2114 286538 2119
rect 286510 240 286538 2086
rect 275100 -480 275212 196
rect 275254 182 275450 210
rect 276052 -480 276164 240
rect 277004 -480 277116 240
rect 277942 196 278068 240
rect 277956 -480 278068 196
rect 278908 -480 279020 240
rect 279860 -480 279972 240
rect 280798 196 280924 240
rect 280812 -480 280924 196
rect 281764 -480 281876 240
rect 282716 -480 282828 240
rect 283654 196 283780 240
rect 283668 -480 283780 196
rect 284620 -480 284732 240
rect 285572 -480 285684 240
rect 286510 196 286636 240
rect 286524 -480 286636 196
rect 287476 -480 287588 240
rect 288428 -480 288540 240
rect 289380 -480 289492 240
rect 290332 -480 290444 240
rect 291284 -480 291396 240
rect 292236 -480 292348 240
<< via2 >>
rect 20398 295246 20426 295274
rect 27566 295246 27594 295274
rect 82838 295638 82866 295666
rect 86926 295638 86954 295666
rect 71806 295414 71834 295442
rect 60774 295358 60802 295386
rect 86086 295358 86114 295386
rect 49742 295302 49770 295330
rect 38710 295246 38738 295274
rect 22918 168406 22946 168434
rect 26950 166726 26978 166754
rect 30982 164206 31010 164234
rect 32326 162526 32354 162554
rect 29638 161854 29666 161882
rect 28294 161798 28322 161826
rect 25606 161742 25634 161770
rect 24262 161686 24290 161714
rect 33670 161294 33698 161322
rect 34062 168406 34090 168434
rect 34734 161686 34762 161714
rect 36078 166726 36106 166754
rect 35014 161686 35042 161714
rect 35406 161742 35434 161770
rect 36358 162078 36386 162106
rect 37422 161854 37450 161882
rect 36750 161798 36778 161826
rect 37702 161798 37730 161826
rect 38094 164206 38122 164234
rect 38766 162526 38794 162554
rect 39046 161854 39074 161882
rect 40110 161686 40138 161714
rect 39438 161294 39466 161322
rect 41734 162134 41762 162162
rect 40390 161294 40418 161322
rect 40782 162078 40810 162106
rect 42126 161854 42154 161882
rect 41454 161798 41482 161826
rect 42798 161294 42826 161322
rect 43078 161294 43106 161322
rect 44142 162134 44170 162162
rect 44422 162078 44450 162106
rect 45486 162078 45514 162106
rect 44814 161294 44842 161322
rect 48174 167230 48202 167258
rect 47502 167174 47530 167202
rect 49798 167230 49826 167258
rect 50190 167734 50218 167762
rect 48454 167174 48482 167202
rect 48846 167174 48874 167202
rect 49518 162974 49546 163002
rect 50862 167678 50890 167706
rect 52206 167566 52234 167594
rect 51142 167174 51170 167202
rect 51534 167174 51562 167202
rect 53830 167734 53858 167762
rect 55174 167678 55202 167706
rect 57862 167566 57890 167594
rect 56518 167174 56546 167202
rect 56910 167006 56938 167034
rect 53550 166894 53578 166922
rect 52486 162974 52514 163002
rect 52878 166726 52906 166754
rect 56238 161686 56266 161714
rect 57582 166950 57610 166978
rect 58254 166838 58282 166866
rect 58926 166782 58954 166810
rect 60270 168630 60298 168658
rect 59206 166726 59234 166754
rect 59598 166726 59626 166754
rect 60550 166894 60578 166922
rect 60942 168574 60970 168602
rect 61614 168406 61642 168434
rect 63238 167006 63266 167034
rect 63406 168518 63434 168546
rect 61894 161686 61922 161714
rect 62286 162078 62314 162106
rect 63406 162078 63434 162106
rect 64414 168462 64442 168490
rect 62958 162022 62986 162050
rect 64582 166950 64610 166978
rect 65926 166838 65954 166866
rect 67270 166782 67298 166810
rect 69958 168630 69986 168658
rect 71302 168574 71330 168602
rect 73990 168518 74018 168546
rect 75334 168462 75362 168490
rect 72646 168406 72674 168434
rect 68614 166726 68642 166754
rect 64414 162022 64442 162050
rect 70966 165046 70994 165074
rect 65646 161966 65674 161994
rect 63630 161910 63658 161938
rect 64302 161854 64330 161882
rect 64974 161798 65002 161826
rect 70966 161966 70994 161994
rect 76678 161910 76706 161938
rect 78022 161854 78050 161882
rect 80710 165046 80738 165074
rect 79366 161798 79394 161826
rect 66318 161742 66346 161770
rect 82054 161742 82082 161770
rect 66990 161686 67018 161714
rect 86086 162078 86114 162106
rect 86478 295246 86506 295274
rect 83398 161686 83426 161714
rect 86926 161350 86954 161378
rect 87038 295414 87066 295442
rect 93646 295414 93674 295442
rect 87038 161294 87066 161322
rect 87150 295302 87178 295330
rect 87822 162078 87850 162106
rect 91854 162078 91882 162106
rect 89838 162022 89866 162050
rect 89166 161350 89194 161378
rect 88494 161294 88522 161322
rect 90510 161798 90538 161826
rect 91182 161686 91210 161714
rect 93646 162078 93674 162106
rect 95326 295526 95354 295554
rect 93758 162022 93786 162050
rect 93870 295246 93898 295274
rect 93198 161742 93226 161770
rect 92526 161294 92554 161322
rect 104790 295526 104818 295554
rect 99526 295470 99554 295498
rect 95326 161798 95354 161826
rect 95438 295358 95466 295386
rect 115822 295470 115850 295498
rect 126854 295414 126882 295442
rect 137886 295358 137914 295386
rect 99638 295302 99666 295330
rect 148918 295302 148946 295330
rect 159950 295246 159978 295274
rect 204190 295414 204218 295442
rect 193158 295358 193186 295386
rect 182126 295302 182154 295330
rect 208726 295302 208754 295330
rect 171094 295246 171122 295274
rect 102606 167286 102634 167314
rect 99638 161742 99666 161770
rect 101934 167174 101962 167202
rect 99526 161686 99554 161714
rect 95438 161294 95466 161322
rect 102942 167174 102970 167202
rect 103278 167342 103306 167370
rect 104286 167286 104314 167314
rect 105294 168014 105322 168042
rect 104622 163758 104650 163786
rect 103950 163422 103978 163450
rect 106638 167902 106666 167930
rect 105630 167342 105658 167370
rect 105966 167342 105994 167370
rect 106974 163422 107002 163450
rect 107310 167846 107338 167874
rect 107982 167790 108010 167818
rect 109662 168014 109690 168042
rect 108318 163758 108346 163786
rect 108654 167734 108682 167762
rect 109326 167678 109354 167706
rect 109998 167622 110026 167650
rect 112350 167902 112378 167930
rect 113694 167846 113722 167874
rect 114702 168630 114730 168658
rect 111006 167342 111034 167370
rect 112014 167566 112042 167594
rect 110670 161854 110698 161882
rect 112686 162526 112714 162554
rect 113358 161798 113386 161826
rect 114030 161742 114058 161770
rect 115038 167790 115066 167818
rect 116046 168574 116074 168602
rect 115374 161686 115402 161714
rect 116382 167734 116410 167762
rect 116718 168518 116746 168546
rect 117390 168462 117418 168490
rect 116774 163758 116802 163786
rect 116774 161854 116802 161882
rect 117726 167678 117754 167706
rect 118062 168406 118090 168434
rect 119070 167622 119098 167650
rect 121758 167566 121786 167594
rect 120414 163758 120442 163786
rect 120078 163422 120106 163450
rect 118734 162078 118762 162106
rect 119406 162022 119434 162050
rect 121422 163366 121450 163394
rect 120750 161910 120778 161938
rect 123102 162526 123130 162554
rect 124110 161966 124138 161994
rect 125566 168686 125594 168714
rect 125566 162078 125594 162106
rect 124446 161798 124474 161826
rect 125454 161854 125482 161882
rect 124782 161630 124810 161658
rect 127134 168630 127162 168658
rect 127470 162638 127498 162666
rect 125790 161742 125818 161770
rect 126126 162526 126154 162554
rect 126798 161798 126826 161826
rect 128142 161742 128170 161770
rect 129822 168574 129850 168602
rect 129934 168630 129962 168658
rect 128478 161686 128506 161714
rect 128814 162582 128842 162610
rect 129486 161686 129514 161714
rect 131166 168518 131194 168546
rect 131614 168574 131642 168602
rect 130830 162862 130858 162890
rect 129934 161630 129962 161658
rect 130158 162134 130186 162162
rect 131502 162806 131530 162834
rect 132286 168518 132314 168546
rect 131614 162526 131642 162554
rect 132174 162750 132202 162778
rect 132510 168462 132538 168490
rect 135198 168686 135226 168714
rect 133854 168406 133882 168434
rect 133966 168462 133994 168490
rect 132286 162638 132314 162666
rect 132846 162694 132874 162722
rect 133518 162638 133546 162666
rect 134974 168406 135002 168434
rect 133966 162582 133994 162610
rect 134190 162582 134218 162610
rect 134862 162526 134890 162554
rect 134974 162134 135002 162162
rect 137886 163422 137914 163450
rect 136542 162022 136570 162050
rect 140574 163366 140602 163394
rect 143262 168630 143290 168658
rect 141918 161966 141946 161994
rect 139230 161910 139258 161938
rect 145950 168574 145978 168602
rect 144606 161854 144634 161882
rect 148638 168518 148666 168546
rect 147294 161798 147322 161826
rect 151326 168462 151354 168490
rect 149982 161742 150010 161770
rect 154014 168406 154042 168434
rect 155358 162862 155386 162890
rect 156702 162806 156730 162834
rect 158046 162750 158074 162778
rect 159390 162694 159418 162722
rect 160734 162638 160762 162666
rect 162078 162582 162106 162610
rect 180558 168574 180586 168602
rect 179886 168518 179914 168546
rect 179214 168462 179242 168490
rect 175854 168406 175882 168434
rect 163422 162526 163450 162554
rect 174510 167566 174538 167594
rect 152670 161686 152698 161714
rect 175182 165886 175210 165914
rect 181006 167566 181034 167594
rect 181230 167230 181258 167258
rect 181566 165886 181594 165914
rect 181902 167174 181930 167202
rect 182126 164598 182154 164626
rect 182574 164598 182602 164626
rect 182686 164598 182714 164626
rect 183246 164598 183274 164626
rect 183806 167230 183834 167258
rect 184366 167174 184394 167202
rect 188846 168574 188874 168602
rect 188286 168518 188314 168546
rect 187726 168406 187754 168434
rect 187950 167230 187978 167258
rect 189406 167230 189434 167258
rect 188622 167174 188650 167202
rect 190526 168462 190554 168490
rect 189966 167174 189994 167202
rect 191646 168630 191674 168658
rect 191086 162022 191114 162050
rect 192206 161966 192234 161994
rect 192766 161910 192794 161938
rect 193886 168518 193914 168546
rect 193326 161854 193354 161882
rect 195006 168462 195034 168490
rect 194446 161798 194474 161826
rect 196126 168406 196154 168434
rect 195566 161742 195594 161770
rect 197246 168574 197274 168602
rect 198366 168686 198394 168714
rect 197806 162638 197834 162666
rect 199486 168742 199514 168770
rect 198926 162526 198954 162554
rect 200046 162470 200074 162498
rect 201166 162862 201194 162890
rect 201726 162806 201754 162834
rect 202062 168630 202090 168658
rect 200606 162414 200634 162442
rect 201166 162638 201194 162666
rect 201166 162078 201194 162106
rect 196686 161686 196714 161714
rect 201390 162022 201418 162050
rect 202286 162750 202314 162778
rect 202846 162694 202874 162722
rect 203406 162638 203434 162666
rect 202454 162526 202482 162554
rect 205534 168742 205562 168770
rect 203966 162526 203994 162554
rect 204750 168518 204778 168546
rect 202454 162022 202482 162050
rect 203294 162470 203322 162498
rect 202734 161966 202762 161994
rect 203294 161966 203322 161994
rect 203518 162414 203546 162442
rect 203406 161910 203434 161938
rect 203518 161910 203546 161938
rect 204078 161854 204106 161882
rect 205422 161798 205450 161826
rect 207046 168686 207074 168714
rect 205534 161798 205562 161826
rect 206094 168462 206122 168490
rect 207886 168574 207914 168602
rect 207438 168406 207466 168434
rect 207158 162022 207186 162050
rect 206766 161742 206794 161770
rect 216398 295414 216426 295442
rect 215110 166726 215138 166754
rect 216286 295358 216314 295386
rect 208726 162582 208754 162610
rect 213486 162862 213514 162890
rect 209454 162078 209482 162106
rect 207886 161294 207914 161322
rect 208110 161686 208138 161714
rect 208782 161294 208810 161322
rect 210126 162022 210154 162050
rect 212142 161966 212170 161994
rect 211470 161798 211498 161826
rect 210798 161742 210826 161770
rect 212814 161910 212842 161938
rect 214158 162806 214186 162834
rect 214830 162750 214858 162778
rect 215502 162694 215530 162722
rect 216174 162638 216202 162666
rect 216286 161742 216314 161770
rect 225582 295302 225610 295330
rect 216398 161686 216426 161714
rect 216510 295246 216538 295274
rect 224686 295078 224714 295106
rect 223566 166726 223594 166754
rect 221550 162582 221578 162610
rect 216510 161294 216538 161322
rect 216846 162526 216874 162554
rect 220878 161294 220906 161322
rect 222222 161742 222250 161770
rect 222894 161686 222922 161714
rect 224238 161294 224266 161322
rect 224686 161294 224714 161322
rect 224910 161294 224938 161322
rect 227206 295358 227234 295386
rect 226142 295078 226170 295106
rect 226254 295246 226282 295274
rect 237174 295358 237202 295386
rect 248206 295302 248234 295330
rect 259238 295246 259266 295274
rect 235662 166278 235690 166306
rect 232974 166222 233002 166250
rect 232302 165942 232330 165970
rect 227206 161294 227234 161322
rect 230286 165886 230314 165914
rect 230958 161686 230986 161714
rect 234990 166166 235018 166194
rect 233646 165830 233674 165858
rect 234318 165774 234346 165802
rect 235886 165886 235914 165914
rect 236334 167734 236362 167762
rect 236558 161686 236586 161714
rect 237006 167622 237034 167650
rect 237230 165942 237258 165970
rect 237678 167566 237706 167594
rect 237902 166222 237930 166250
rect 238350 167678 238378 167706
rect 238574 165830 238602 165858
rect 239022 167958 239050 167986
rect 239246 165774 239274 165802
rect 239694 167174 239722 167202
rect 239918 166166 239946 166194
rect 240366 167902 240394 167930
rect 240590 166278 240618 166306
rect 241038 167846 241066 167874
rect 241262 167734 241290 167762
rect 241934 167622 241962 167650
rect 243950 167958 243978 167986
rect 243278 167678 243306 167706
rect 242606 167566 242634 167594
rect 245294 167902 245322 167930
rect 245966 167846 245994 167874
rect 244622 167174 244650 167202
rect 247982 165998 248010 166026
rect 248654 165886 248682 165914
rect 247310 164318 247338 164346
rect 246638 164206 246666 164234
rect 249998 164262 250026 164290
rect 249326 163422 249354 163450
rect 251342 165942 251370 165970
rect 250670 163366 250698 163394
rect 253358 165046 253386 165074
rect 253806 164318 253834 164346
rect 252686 162582 252714 162610
rect 253134 164206 253162 164234
rect 252014 162526 252042 162554
rect 254702 168406 254730 168434
rect 261198 168406 261226 168434
rect 254030 163478 254058 163506
rect 254478 165998 254506 166026
rect 257838 165942 257866 165970
rect 255150 165886 255178 165914
rect 256494 164262 256522 164290
rect 255822 163422 255850 163450
rect 257166 163366 257194 163394
rect 259854 165046 259882 165074
rect 259182 162582 259210 162610
rect 258510 162526 258538 162554
rect 260526 163478 260554 163506
rect 269710 159334 269738 159362
rect 273406 295246 273434 295274
rect 281302 295246 281330 295274
rect 273406 158550 273434 158578
rect 292334 158102 292362 158130
rect 20398 157766 20426 157794
rect 16534 157206 16562 157234
rect 5502 156646 5530 156674
rect 277606 137494 277634 137522
rect 275422 135646 275450 135674
rect 272118 135254 272146 135282
rect 33950 129038 33978 129066
rect 16814 128982 16842 129010
rect 24430 107086 24458 107114
rect 22526 106358 22554 106386
rect 18718 106302 18746 106330
rect 20622 106246 20650 106274
rect 30142 106582 30170 106610
rect 28238 106470 28266 106498
rect 26334 106414 26362 106442
rect 32046 106526 32074 106554
rect 35070 128982 35098 129010
rect 34846 128926 34874 128954
rect 34846 106302 34874 106330
rect 35854 107142 35882 107170
rect 37366 128982 37394 129010
rect 37366 106582 37394 106610
rect 39102 106414 39130 106442
rect 39662 106582 39690 106610
rect 37758 106358 37786 106386
rect 37086 106246 37114 106274
rect 37758 106246 37786 106274
rect 41790 129038 41818 129066
rect 41118 106526 41146 106554
rect 41566 107198 41594 107226
rect 39774 106470 39802 106498
rect 43134 106246 43162 106274
rect 43470 106638 43498 106666
rect 45150 106638 45178 106666
rect 43806 106582 43834 106610
rect 47838 128870 47866 128898
rect 48286 128870 48314 128898
rect 47166 106638 47194 106666
rect 47278 107254 47306 107282
rect 49182 128870 49210 128898
rect 48286 106582 48314 106610
rect 49182 106638 49210 106666
rect 49966 128870 49994 128898
rect 51198 128534 51226 128562
rect 51646 128534 51674 128562
rect 49966 106358 49994 106386
rect 51086 106582 51114 106610
rect 49854 106302 49882 106330
rect 51870 106582 51898 106610
rect 52990 107310 53018 107338
rect 51646 106246 51674 106274
rect 53886 129038 53914 129066
rect 55902 129094 55930 129122
rect 57246 107366 57274 107394
rect 55230 106526 55258 106554
rect 57918 106470 57946 106498
rect 58702 107422 58730 107450
rect 53214 106414 53242 106442
rect 54894 106358 54922 106386
rect 56798 106302 56826 106330
rect 59262 106358 59290 106386
rect 59934 106302 59962 106330
rect 60606 106246 60634 106274
rect 61950 129206 61978 129234
rect 66990 129206 67018 129234
rect 66766 129150 66794 129178
rect 64414 106638 64442 106666
rect 61278 106246 61306 106274
rect 62510 106582 62538 106610
rect 66766 106638 66794 106666
rect 66878 129038 66906 129066
rect 66878 106638 66906 106666
rect 66318 106414 66346 106442
rect 68446 129094 68474 129122
rect 66990 106414 67018 106442
rect 68222 106638 68250 106666
rect 68446 106582 68474 106610
rect 70126 129038 70154 129066
rect 70686 128926 70714 128954
rect 72030 128982 72058 129010
rect 76062 129150 76090 129178
rect 76734 129038 76762 129066
rect 75390 107422 75418 107450
rect 75838 128870 75866 128898
rect 74718 107310 74746 107338
rect 74046 107254 74074 107282
rect 73374 107198 73402 107226
rect 72702 107142 72730 107170
rect 71358 107086 71386 107114
rect 73934 106582 73962 106610
rect 72030 106526 72058 106554
rect 77406 128870 77434 128898
rect 77742 107366 77770 107394
rect 78078 106638 78106 106666
rect 82782 127246 82810 127274
rect 84798 127302 84826 127330
rect 83454 126574 83482 126602
rect 86142 128926 86170 128954
rect 86814 127358 86842 127386
rect 90174 128982 90202 129010
rect 89502 128086 89530 128114
rect 88830 127414 88858 127442
rect 91518 129206 91546 129234
rect 90846 126742 90874 126770
rect 94206 129038 94234 129066
rect 93534 128142 93562 128170
rect 92862 127470 92890 127498
rect 92190 126630 92218 126658
rect 88158 126518 88186 126546
rect 87486 126462 87514 126490
rect 85470 126406 85498 126434
rect 95550 129262 95578 129290
rect 97566 129318 97594 129346
rect 96894 129150 96922 129178
rect 98238 129094 98266 129122
rect 98910 128366 98938 128394
rect 99134 129206 99162 129234
rect 99582 128198 99610 128226
rect 99134 127526 99162 127554
rect 100926 129206 100954 129234
rect 101598 128254 101626 128282
rect 100254 126798 100282 126826
rect 102046 127246 102074 127274
rect 96222 126686 96250 126714
rect 94878 126350 94906 126378
rect 102886 129318 102914 129346
rect 102438 129262 102466 129290
rect 102886 127638 102914 127666
rect 102438 127582 102466 127610
rect 102270 127246 102298 127274
rect 102494 127302 102522 127330
rect 102270 126574 102298 126602
rect 102942 127190 102970 127218
rect 103166 127358 103194 127386
rect 103614 126574 103642 126602
rect 103838 127414 103866 127442
rect 104958 126854 104986 126882
rect 105182 127470 105210 127498
rect 104286 126294 104314 126322
rect 104510 126742 104538 126770
rect 106302 128310 106330 128338
rect 106526 129150 106554 129178
rect 105630 127302 105658 127330
rect 105854 126350 105882 126378
rect 106806 128982 106834 129010
rect 106806 128478 106834 128506
rect 106974 126126 107002 126154
rect 107198 128366 107226 128394
rect 107646 127358 107674 127386
rect 107870 129206 107898 129234
rect 108150 128926 108178 128954
rect 108094 126406 108122 126434
rect 108318 127414 108346 127442
rect 108542 127190 108570 127218
rect 108990 126742 109018 126770
rect 109046 129038 109074 129066
rect 108990 126518 109018 126546
rect 108766 126462 108794 126490
rect 109494 128478 109522 128506
rect 109438 128086 109466 128114
rect 109046 126462 109074 126490
rect 109214 126854 109242 126882
rect 109662 127470 109690 127498
rect 110054 129094 110082 129122
rect 109886 126126 109914 126154
rect 110782 128142 110810 128170
rect 110054 126126 110082 126154
rect 110110 127526 110138 127554
rect 110334 126630 110362 126658
rect 110390 126406 110418 126434
rect 110558 126742 110586 126770
rect 111006 126462 111034 126490
rect 112350 128646 112378 128674
rect 112574 128870 112602 128898
rect 111678 128142 111706 128170
rect 112126 127638 112154 127666
rect 111454 127582 111482 127610
rect 111902 126854 111930 126882
rect 111678 126350 111706 126378
rect 112350 126126 112378 126154
rect 112798 128198 112826 128226
rect 113022 126854 113050 126882
rect 113246 128590 113274 128618
rect 112854 126798 112882 126826
rect 113470 128254 113498 128282
rect 113694 127246 113722 127274
rect 113750 126798 113778 126826
rect 114142 126574 114170 126602
rect 113918 126462 113946 126490
rect 114366 126574 114394 126602
rect 114590 129038 114618 129066
rect 114366 126294 114394 126322
rect 115038 128870 115066 128898
rect 115262 128982 115290 129010
rect 115038 128310 115066 128338
rect 114814 127302 114842 127330
rect 115542 127414 115570 127442
rect 115486 127358 115514 127386
rect 115710 126630 115738 126658
rect 115934 128926 115962 128954
rect 116158 127470 116186 127498
rect 116886 128646 116914 128674
rect 116830 128142 116858 128170
rect 116382 126518 116410 126546
rect 116606 128086 116634 128114
rect 116382 126406 116410 126434
rect 117726 128870 117754 128898
rect 118398 128814 118426 128842
rect 118622 129262 118650 129290
rect 117054 128590 117082 128618
rect 117502 126798 117530 126826
rect 117278 126406 117306 126434
rect 118174 126630 118202 126658
rect 117726 126574 117754 126602
rect 117950 126574 117978 126602
rect 118398 126518 118426 126546
rect 118846 128870 118874 128898
rect 119294 129150 119322 129178
rect 119014 126462 119042 126490
rect 119070 128814 119098 128842
rect 120190 126910 120218 126938
rect 119742 126854 119770 126882
rect 119966 126686 119994 126714
rect 121086 129038 121114 129066
rect 121310 129206 121338 129234
rect 120638 128870 120666 128898
rect 120414 126854 120442 126882
rect 120526 128534 120554 128562
rect 121758 126910 121786 126938
rect 121982 129094 122010 129122
rect 123102 128982 123130 129010
rect 123774 128926 123802 128954
rect 122430 128534 122458 128562
rect 124446 128086 124474 128114
rect 124670 129318 124698 129346
rect 122654 126630 122682 126658
rect 123326 126518 123354 126546
rect 123998 126462 124026 126490
rect 126462 129262 126490 129290
rect 126686 129262 126714 129290
rect 125790 126574 125818 126602
rect 126014 129038 126042 129066
rect 125118 126406 125146 126434
rect 125342 126406 125370 126434
rect 127134 129150 127162 129178
rect 127358 128982 127386 129010
rect 129150 129206 129178 129234
rect 129822 129094 129850 129122
rect 128478 128870 128506 128898
rect 127806 126686 127834 126714
rect 130494 126630 130522 126658
rect 131166 126574 131194 126602
rect 132510 129318 132538 129346
rect 131838 126462 131866 126490
rect 132286 128926 132314 128954
rect 78750 106526 78778 106554
rect 81550 106638 81578 106666
rect 79646 106470 79674 106498
rect 87262 106526 87290 106554
rect 83454 106358 83482 106386
rect 85358 106302 85386 106330
rect 91070 106414 91098 106442
rect 89166 106246 89194 106274
rect 19278 75334 19306 75362
rect 19278 75110 19306 75138
rect 18886 74718 18914 74746
rect 16142 73710 16170 73738
rect 14294 73654 14322 73682
rect 13286 73598 13314 73626
rect 10430 73542 10458 73570
rect 9478 73486 9506 73514
rect 7574 7126 7602 7154
rect 6678 2142 6706 2170
rect 5782 2086 5810 2114
rect 8638 2926 8666 2954
rect 12446 2982 12474 3010
rect 11494 2198 11522 2226
rect 15302 3038 15330 3066
rect 18494 73094 18522 73122
rect 18158 3150 18186 3178
rect 17206 3094 17234 3122
rect 18494 2142 18522 2170
rect 19278 73094 19306 73122
rect 19950 7126 19978 7154
rect 21966 73542 21994 73570
rect 21294 73486 21322 73514
rect 21854 73486 21882 73514
rect 20622 2926 20650 2954
rect 20958 2366 20986 2394
rect 20062 2142 20090 2170
rect 18886 2086 18914 2114
rect 19110 2086 19138 2114
rect 24654 73654 24682 73682
rect 23982 73598 24010 73626
rect 24766 73598 24794 73626
rect 23310 2982 23338 3010
rect 23926 73542 23954 73570
rect 22638 2198 22666 2226
rect 22918 2142 22946 2170
rect 24038 73150 24066 73178
rect 24038 2254 24066 2282
rect 23926 2142 23954 2170
rect 23870 2030 23898 2058
rect 24878 73094 24906 73122
rect 25998 73710 26026 73738
rect 26446 73766 26474 73794
rect 25326 3038 25354 3066
rect 24878 2366 24906 2394
rect 24766 2030 24794 2058
rect 24822 2198 24850 2226
rect 27342 3150 27370 3178
rect 26670 3094 26698 3122
rect 27678 2254 27706 2282
rect 26446 2198 26474 2226
rect 26726 2198 26754 2226
rect 25774 2142 25802 2170
rect 28014 2086 28042 2114
rect 28574 73654 28602 73682
rect 28686 73150 28714 73178
rect 29358 73094 29386 73122
rect 29470 73710 29498 73738
rect 32046 73766 32074 73794
rect 31374 73598 31402 73626
rect 30702 73542 30730 73570
rect 30030 73486 30058 73514
rect 30422 73486 30450 73514
rect 32438 2310 32466 2338
rect 31486 2086 31514 2114
rect 35406 73710 35434 73738
rect 34734 73654 34762 73682
rect 36078 73486 36106 73514
rect 34062 2366 34090 2394
rect 34846 73094 34874 73122
rect 33334 2198 33362 2226
rect 33390 2254 33418 2282
rect 32718 2142 32746 2170
rect 34342 2086 34370 2114
rect 36246 2422 36274 2450
rect 34846 2086 34874 2114
rect 35238 2086 35266 2114
rect 36750 2142 36778 2170
rect 37198 2478 37226 2506
rect 37422 2310 37450 2338
rect 38766 73094 38794 73122
rect 38990 73486 39018 73514
rect 38094 2254 38122 2282
rect 38150 2310 38178 2338
rect 40782 2478 40810 2506
rect 40110 2422 40138 2450
rect 42126 73486 42154 73514
rect 41454 2310 41482 2338
rect 41846 73150 41874 73178
rect 41006 2142 41034 2170
rect 39438 2086 39466 2114
rect 40054 2086 40082 2114
rect 44142 73150 44170 73178
rect 43470 2142 43498 2170
rect 43750 73094 43778 73122
rect 42798 2086 42826 2114
rect 42910 2086 42938 2114
rect 45486 73094 45514 73122
rect 44758 2086 44786 2114
rect 44814 2422 44842 2450
rect 46158 2422 46186 2450
rect 45766 2142 45794 2170
rect 46830 2142 46858 2170
rect 46718 2086 46746 2114
rect 47502 2086 47530 2114
rect 47670 2086 47698 2114
rect 48174 2086 48202 2114
rect 52206 73150 52234 73178
rect 51534 73094 51562 73122
rect 52318 73094 52346 73122
rect 52878 73094 52906 73122
rect 53270 73150 53298 73178
rect 54222 73262 54250 73290
rect 54894 73206 54922 73234
rect 53550 73150 53578 73178
rect 55174 73150 55202 73178
rect 54166 73094 54194 73122
rect 55566 2478 55594 2506
rect 56126 73262 56154 73290
rect 56910 73542 56938 73570
rect 56238 2198 56266 2226
rect 57134 73206 57162 73234
rect 57582 2086 57610 2114
rect 58030 2478 58058 2506
rect 58926 73094 58954 73122
rect 59598 2478 59626 2506
rect 59934 73542 59962 73570
rect 58254 2030 58282 2058
rect 58982 2198 59010 2226
rect 60942 2254 60970 2282
rect 60270 2198 60298 2226
rect 62286 73598 62314 73626
rect 62958 73486 62986 73514
rect 61614 2142 61642 2170
rect 62790 73094 62818 73122
rect 60886 2086 60914 2114
rect 61838 2030 61866 2058
rect 64974 73206 65002 73234
rect 65198 73598 65226 73626
rect 64302 73094 64330 73122
rect 65086 73094 65114 73122
rect 63630 2030 63658 2058
rect 63742 2478 63770 2506
rect 65086 2422 65114 2450
rect 64694 2198 64722 2226
rect 66990 73598 67018 73626
rect 66318 73150 66346 73178
rect 65646 73094 65674 73122
rect 66766 73094 66794 73122
rect 65198 2086 65226 2114
rect 65646 2254 65674 2282
rect 66598 2142 66626 2170
rect 67662 2254 67690 2282
rect 67774 73486 67802 73514
rect 66766 2142 66794 2170
rect 67550 2086 67578 2114
rect 68334 73486 68362 73514
rect 68446 73150 68474 73178
rect 69006 73094 69034 73122
rect 69286 73206 69314 73234
rect 68446 2310 68474 2338
rect 67774 2086 67802 2114
rect 68502 2086 68530 2114
rect 69678 3206 69706 3234
rect 70350 3150 70378 3178
rect 70966 73598 70994 73626
rect 70406 2422 70434 2450
rect 69286 2030 69314 2058
rect 69454 2086 69482 2114
rect 71022 73150 71050 73178
rect 71694 3094 71722 3122
rect 72366 3038 72394 3066
rect 72646 73486 72674 73514
rect 72646 2422 72674 2450
rect 72758 73094 72786 73122
rect 73038 73094 73066 73122
rect 73486 73150 73514 73178
rect 72758 2198 72786 2226
rect 73262 2310 73290 2338
rect 70966 2086 70994 2114
rect 72310 2142 72338 2170
rect 71414 2030 71442 2058
rect 74382 73542 74410 73570
rect 73710 2982 73738 3010
rect 73486 2310 73514 2338
rect 74214 2086 74242 2114
rect 75166 73094 75194 73122
rect 75054 2086 75082 2114
rect 75166 2254 75194 2282
rect 75726 3318 75754 3346
rect 77070 73598 77098 73626
rect 77742 3262 77770 3290
rect 76398 2926 76426 2954
rect 78022 3206 78050 3234
rect 75222 2142 75250 2170
rect 76118 2422 76146 2450
rect 77070 2198 77098 2226
rect 79086 73710 79114 73738
rect 79758 73094 79786 73122
rect 80206 73094 80234 73122
rect 80206 3206 80234 3234
rect 78414 2198 78442 2226
rect 78974 3150 79002 3178
rect 81102 73486 81130 73514
rect 80430 3150 80458 3178
rect 80878 3094 80906 3122
rect 79926 2310 79954 2338
rect 82446 73822 82474 73850
rect 81774 3094 81802 3122
rect 81830 3038 81858 3066
rect 82782 2142 82810 2170
rect 84462 73878 84490 73906
rect 83790 3038 83818 3066
rect 84686 73542 84714 73570
rect 83118 2142 83146 2170
rect 83734 2982 83762 3010
rect 85134 73542 85162 73570
rect 85806 2982 85834 3010
rect 85694 2086 85722 2114
rect 87150 73654 87178 73682
rect 87766 73598 87794 73626
rect 86478 2086 86506 2114
rect 86590 3318 86618 3346
rect 87542 2926 87570 2954
rect 88494 73766 88522 73794
rect 87822 2926 87850 2954
rect 88606 73710 88634 73738
rect 90286 73878 90314 73906
rect 89166 73598 89194 73626
rect 89502 73822 89530 73850
rect 88606 2534 88634 2562
rect 89446 3262 89474 3290
rect 87766 2030 87794 2058
rect 88494 2030 88522 2058
rect 89502 2310 89530 2338
rect 96166 73766 96194 73794
rect 93646 73486 93674 73514
rect 92302 3206 92330 3234
rect 90286 2254 90314 2282
rect 91350 2534 91378 2562
rect 90398 2198 90426 2226
rect 93254 3150 93282 3178
rect 97846 73654 97874 73682
rect 96278 73542 96306 73570
rect 95158 3094 95186 3122
rect 93646 2142 93674 2170
rect 94206 2142 94234 2170
rect 96110 2310 96138 2338
rect 96278 2366 96306 2394
rect 96222 2310 96250 2338
rect 97230 2310 97258 2338
rect 99526 73598 99554 73626
rect 97846 2310 97874 2338
rect 98014 3038 98042 3066
rect 97230 2198 97258 2226
rect 97062 2142 97090 2170
rect 98966 2254 98994 2282
rect 100870 2982 100898 3010
rect 99526 2142 99554 2170
rect 99974 2366 100002 2394
rect 103726 2926 103754 2954
rect 102774 2310 102802 2338
rect 101822 2086 101850 2114
rect 104678 2198 104706 2226
rect 105630 2142 105658 2170
rect 129542 2086 129570 2114
rect 134526 129262 134554 129290
rect 133854 129038 133882 129066
rect 135198 128982 135226 129010
rect 137998 128982 138026 129010
rect 133182 126406 133210 126434
rect 135198 2142 135226 2170
rect 143262 128926 143290 128954
rect 142590 2086 142618 2114
rect 143822 2478 143850 2506
rect 140966 2030 140994 2058
rect 144606 128982 144634 129010
rect 143934 2142 143962 2170
rect 145950 2478 145978 2506
rect 145278 2030 145306 2058
rect 148638 128982 148666 129010
rect 149982 128926 150010 128954
rect 149310 2926 149338 2954
rect 147966 2422 147994 2450
rect 150654 2254 150682 2282
rect 151326 2198 151354 2226
rect 151998 2142 152026 2170
rect 152278 2422 152306 2450
rect 147294 2086 147322 2114
rect 149422 2086 149450 2114
rect 172102 129094 172130 129122
rect 170982 129038 171010 129066
rect 152670 2086 152698 2114
rect 155134 128982 155162 129010
rect 169862 128982 169890 129010
rect 159166 128926 159194 128954
rect 157990 2926 158018 2954
rect 163142 128926 163170 128954
rect 168742 126518 168770 126546
rect 167622 126462 167650 126490
rect 166502 126406 166530 126434
rect 173502 128926 173530 128954
rect 174342 128926 174370 128954
rect 173222 126574 173250 126602
rect 175462 128086 175490 128114
rect 176190 126462 176218 126490
rect 176582 126798 176610 126826
rect 175518 126406 175546 126434
rect 178878 129094 178906 129122
rect 178206 129038 178234 129066
rect 178822 129038 178850 129066
rect 177534 128982 177562 129010
rect 176862 126518 176890 126546
rect 177702 128534 177730 128562
rect 179550 126574 179578 126602
rect 179942 129094 179970 129122
rect 180222 128926 180250 128954
rect 180894 128086 180922 128114
rect 181062 128870 181090 128898
rect 181566 126798 181594 126826
rect 182182 128926 182210 128954
rect 183582 129094 183610 129122
rect 182910 129038 182938 129066
rect 184926 128926 184954 128954
rect 184254 128870 184282 128898
rect 184422 128870 184450 128898
rect 182238 128534 182266 128562
rect 183302 128814 183330 128842
rect 186270 128870 186298 128898
rect 185598 128814 185626 128842
rect 185542 128534 185570 128562
rect 186942 128534 186970 128562
rect 186662 126854 186690 126882
rect 187614 126854 187642 126882
rect 190302 128870 190330 128898
rect 190974 128814 191002 128842
rect 191142 128870 191170 128898
rect 191646 126798 191674 126826
rect 192262 128814 192290 128842
rect 192318 126406 192346 126434
rect 192990 126238 193018 126266
rect 193382 126798 193410 126826
rect 193662 126182 193690 126210
rect 195678 129038 195706 129066
rect 196350 128982 196378 129010
rect 197022 128926 197050 128954
rect 197694 128142 197722 128170
rect 198366 128086 198394 128114
rect 195006 126742 195034 126770
rect 198982 126742 199010 126770
rect 194334 126126 194362 126154
rect 194502 126406 194530 126434
rect 195622 126238 195650 126266
rect 196742 126182 196770 126210
rect 197862 126126 197890 126154
rect 199710 127302 199738 127330
rect 200102 129038 200130 129066
rect 199038 126686 199066 126714
rect 200382 126630 200410 126658
rect 201054 126574 201082 126602
rect 201222 128982 201250 129010
rect 201726 127246 201754 127274
rect 202342 128926 202370 128954
rect 203742 129094 203770 129122
rect 204414 128926 204442 128954
rect 203070 127526 203098 127554
rect 203462 128142 203490 128170
rect 202398 126518 202426 126546
rect 204582 128086 204610 128114
rect 205086 126462 205114 126490
rect 205702 126686 205730 126714
rect 205758 126406 205786 126434
rect 206430 126350 206458 126378
rect 206822 127302 206850 127330
rect 207774 127470 207802 127498
rect 208446 127414 208474 127442
rect 209118 127358 209146 127386
rect 210462 129038 210490 129066
rect 209790 127302 209818 127330
rect 207102 126798 207130 126826
rect 210182 127246 210210 127274
rect 207942 126630 207970 126658
rect 209062 126574 209090 126602
rect 211806 128982 211834 129010
rect 212478 128086 212506 128114
rect 211134 127246 211162 127274
rect 212422 127526 212450 127554
rect 211302 126518 211330 126546
rect 213150 126742 213178 126770
rect 213542 129094 213570 129122
rect 213822 126686 213850 126714
rect 214494 126630 214522 126658
rect 214662 128926 214690 128954
rect 215166 126574 215194 126602
rect 215838 126518 215866 126546
rect 215782 126462 215810 126490
rect 216510 126462 216538 126490
rect 216902 126406 216930 126434
rect 223230 129206 223258 129234
rect 222558 129094 222586 129122
rect 217854 128926 217882 128954
rect 224574 129150 224602 129178
rect 223902 128534 223930 128562
rect 224742 129038 224770 129066
rect 220262 127470 220290 127498
rect 217182 126406 217210 126434
rect 219142 126798 219170 126826
rect 218022 126350 218050 126378
rect 221382 127414 221410 127442
rect 222502 127358 222530 127386
rect 223622 127302 223650 127330
rect 225246 127526 225274 127554
rect 225862 127246 225890 127274
rect 226590 127470 226618 127498
rect 226982 128982 227010 129010
rect 225918 126798 225946 126826
rect 227262 127414 227290 127442
rect 228494 128534 228522 128562
rect 227934 127358 227962 127386
rect 228102 128086 228130 128114
rect 228606 127302 228634 127330
rect 229950 128310 229978 128338
rect 230622 128254 230650 128282
rect 230958 129206 230986 129234
rect 229278 127246 229306 127274
rect 228494 126350 228522 126378
rect 229222 126742 229250 126770
rect 230342 126686 230370 126714
rect 231294 128198 231322 128226
rect 231798 129094 231826 129122
rect 230958 126238 230986 126266
rect 231462 126630 231490 126658
rect 231966 128142 231994 128170
rect 232246 129150 232274 129178
rect 231798 126630 231826 126658
rect 233310 129262 233338 129290
rect 233982 129206 234010 129234
rect 234654 129094 234682 129122
rect 232638 128982 232666 129010
rect 233814 128926 233842 128954
rect 232246 126294 232274 126322
rect 232582 126574 232610 126602
rect 233702 126518 233730 126546
rect 236670 129318 236698 129346
rect 235998 129038 236026 129066
rect 237342 128926 237370 128954
rect 235326 128086 235354 128114
rect 238014 126742 238042 126770
rect 238686 126686 238714 126714
rect 238182 126630 238210 126658
rect 233814 126182 233842 126210
rect 234822 126462 234850 126490
rect 235942 126406 235970 126434
rect 237062 126182 237090 126210
rect 239414 128982 239442 129010
rect 240030 128982 240058 129010
rect 239414 127582 239442 127610
rect 239358 126630 239386 126658
rect 241374 129150 241402 129178
rect 240702 126574 240730 126602
rect 242046 126518 242074 126546
rect 242718 129262 242746 129290
rect 242718 127638 242746 127666
rect 242606 126462 242634 126490
rect 242662 127526 242690 127554
rect 240422 126350 240450 126378
rect 239302 126238 239330 126266
rect 241542 126294 241570 126322
rect 245014 129318 245042 129346
rect 243558 129206 243586 129234
rect 243558 127526 243586 127554
rect 244902 127470 244930 127498
rect 243390 126406 243418 126434
rect 243782 126798 243810 126826
rect 251566 129150 251594 129178
rect 245014 127470 245042 127498
rect 250502 128478 250530 128506
rect 246022 127414 246050 127442
rect 247142 127358 247170 127386
rect 248262 127302 248290 127330
rect 249382 127246 249410 127274
rect 258342 129094 258370 129122
rect 251566 128254 251594 128282
rect 251622 128422 251650 128450
rect 252742 128142 252770 128170
rect 253862 128030 253890 128058
rect 256102 127638 256130 127666
rect 254982 127582 255010 127610
rect 257222 127526 257250 127554
rect 260582 129038 260610 129066
rect 259462 128086 259490 128114
rect 265398 128982 265426 129010
rect 262822 128926 262850 128954
rect 261702 127470 261730 127498
rect 263942 126742 263970 126770
rect 265062 126686 265090 126714
rect 269542 128254 269570 128282
rect 265398 126182 265426 126210
rect 266182 126630 266210 126658
rect 268422 126574 268450 126602
rect 267302 126182 267330 126210
rect 270662 126518 270690 126546
rect 271782 126462 271810 126490
rect 272902 126406 272930 126434
rect 272118 124782 272146 124810
rect 269374 7126 269402 7154
rect 260806 6398 260834 6426
rect 249382 6342 249410 6370
rect 243670 6286 243698 6314
rect 163702 2254 163730 2282
rect 159166 2030 159194 2058
rect 160846 2030 160874 2058
rect 166558 2198 166586 2226
rect 169414 2142 169442 2170
rect 172270 2086 172298 2114
rect 246638 3766 246666 3794
rect 252350 4606 252378 4634
rect 255206 3822 255234 3850
rect 258062 2926 258090 2954
rect 266630 3038 266658 3066
rect 263718 2982 263746 3010
rect 272342 2086 272370 2114
rect 276430 134358 276458 134386
rect 276374 133910 276402 133938
rect 275590 133014 275618 133042
rect 275646 132566 275674 132594
rect 275646 3822 275674 3850
rect 277214 131670 277242 131698
rect 276430 3038 276458 3066
rect 276486 124782 276514 124810
rect 276374 2982 276402 3010
rect 275590 2926 275618 2954
rect 277214 6342 277242 6370
rect 276486 2086 276514 2114
rect 277718 137046 277746 137074
rect 277830 136598 277858 136626
rect 277830 2478 277858 2506
rect 277942 136150 277970 136178
rect 277718 2142 277746 2170
rect 277606 2086 277634 2114
rect 278166 134806 278194 134834
rect 278054 132118 278082 132146
rect 278054 4606 278082 4634
rect 278110 131222 278138 131250
rect 278166 7126 278194 7154
rect 278222 133462 278250 133490
rect 278222 6398 278250 6426
rect 278278 130774 278306 130802
rect 278278 6286 278306 6314
rect 278110 3766 278138 3794
rect 280798 2478 280826 2506
rect 283654 2142 283682 2170
rect 286510 2086 286538 2114
<< metal3 >>
rect 82833 295638 82838 295666
rect 82866 295638 86926 295666
rect 86954 295638 86959 295666
rect 95321 295526 95326 295554
rect 95354 295526 104790 295554
rect 104818 295526 104823 295554
rect 99521 295470 99526 295498
rect 99554 295470 115822 295498
rect 115850 295470 115855 295498
rect 71801 295414 71806 295442
rect 71834 295414 87038 295442
rect 87066 295414 87071 295442
rect 93641 295414 93646 295442
rect 93674 295414 126854 295442
rect 126882 295414 126887 295442
rect 204185 295414 204190 295442
rect 204218 295414 216398 295442
rect 216426 295414 216431 295442
rect 60769 295358 60774 295386
rect 60802 295358 86086 295386
rect 86114 295358 86119 295386
rect 95433 295358 95438 295386
rect 95466 295358 137886 295386
rect 137914 295358 137919 295386
rect 193153 295358 193158 295386
rect 193186 295358 216286 295386
rect 216314 295358 216319 295386
rect 227201 295358 227206 295386
rect 227234 295358 237174 295386
rect 237202 295358 237207 295386
rect 49737 295302 49742 295330
rect 49770 295302 87150 295330
rect 87178 295302 87183 295330
rect 99633 295302 99638 295330
rect 99666 295302 148918 295330
rect 148946 295302 148951 295330
rect 182121 295302 182126 295330
rect 182154 295302 208726 295330
rect 208754 295302 208759 295330
rect 225577 295302 225582 295330
rect 225610 295302 248206 295330
rect 248234 295302 248239 295330
rect 20393 295246 20398 295274
rect 20426 295246 27566 295274
rect 27594 295246 27599 295274
rect 38705 295246 38710 295274
rect 38738 295246 86478 295274
rect 86506 295246 86511 295274
rect 93865 295246 93870 295274
rect 93898 295246 159950 295274
rect 159978 295246 159983 295274
rect 171089 295246 171094 295274
rect 171122 295246 216510 295274
rect 216538 295246 216543 295274
rect 226249 295246 226254 295274
rect 226282 295246 259238 295274
rect 259266 295246 259271 295274
rect 273401 295246 273406 295274
rect 273434 295246 281302 295274
rect 281330 295246 281335 295274
rect 224681 295078 224686 295106
rect 224714 295078 226142 295106
rect 226170 295078 226175 295106
rect 297780 294322 298500 294420
rect 275921 294294 275926 294322
rect 275954 294308 298500 294322
rect 275954 294294 297836 294308
rect -480 293594 240 293692
rect -480 293580 3766 293594
rect 196 293566 3766 293580
rect 3794 293566 3799 293594
rect 297780 287714 298500 287812
rect 271721 287686 271726 287714
rect 271754 287700 298500 287714
rect 271754 287686 297836 287700
rect -480 286538 240 286636
rect -480 286524 2086 286538
rect 196 286510 2086 286524
rect 2114 286510 2119 286538
rect 297780 281106 298500 281204
rect 295241 281078 295246 281106
rect 295274 281092 298500 281106
rect 295274 281078 297836 281092
rect -480 279482 240 279580
rect -480 279468 5446 279482
rect 196 279454 5446 279468
rect 5474 279454 5479 279482
rect 297780 274498 298500 274596
rect 275081 274470 275086 274498
rect 275114 274484 298500 274498
rect 275114 274470 297836 274484
rect -480 272426 240 272524
rect -480 272412 3094 272426
rect 196 272398 3094 272412
rect 3122 272398 3127 272426
rect 297780 267890 298500 267988
rect 278441 267862 278446 267890
rect 278474 267876 298500 267890
rect 278474 267862 297836 267876
rect -480 265370 240 265468
rect -480 265356 2142 265370
rect 196 265342 2142 265356
rect 2170 265342 2175 265370
rect 297780 261282 298500 261380
rect 295297 261254 295302 261282
rect 295330 261268 298500 261282
rect 295330 261254 297836 261268
rect -480 258314 240 258412
rect -480 258300 5502 258314
rect 196 258286 5502 258300
rect 5530 258286 5535 258314
rect 297780 254674 298500 254772
rect 272561 254646 272566 254674
rect 272594 254660 298500 254674
rect 272594 254646 297836 254660
rect -480 251258 240 251356
rect -480 251244 3822 251258
rect 196 251230 3822 251244
rect 3850 251230 3855 251258
rect 297780 248066 298500 248164
rect 272617 248038 272622 248066
rect 272650 248052 298500 248066
rect 272650 248038 297836 248052
rect -480 244202 240 244300
rect -480 244188 2198 244202
rect 196 244174 2198 244188
rect 2226 244174 2231 244202
rect 297780 241458 298500 241556
rect 295353 241430 295358 241458
rect 295386 241444 298500 241458
rect 295386 241430 297836 241444
rect -480 237146 240 237244
rect -480 237132 5558 237146
rect 196 237118 5558 237132
rect 5586 237118 5591 237146
rect 297780 234850 298500 234948
rect 273401 234822 273406 234850
rect 273434 234836 298500 234850
rect 273434 234822 297836 234836
rect -480 230090 240 230188
rect -480 230076 3878 230090
rect 196 230062 3878 230076
rect 3906 230062 3911 230090
rect 297780 228242 298500 228340
rect 277601 228214 277606 228242
rect 277634 228228 298500 228242
rect 277634 228214 297836 228228
rect -480 223034 240 223132
rect -480 223020 2254 223034
rect 196 223006 2254 223020
rect 2282 223006 2287 223034
rect 297780 221634 298500 221732
rect 295409 221606 295414 221634
rect 295442 221620 298500 221634
rect 295442 221606 297836 221620
rect -480 215978 240 216076
rect -480 215964 5614 215978
rect 196 215950 5614 215964
rect 5642 215950 5647 215978
rect 297780 215082 298500 215124
rect 272673 215054 272678 215082
rect 272706 215054 298500 215082
rect 297780 215012 298500 215054
rect -480 208922 240 209020
rect -480 208908 3934 208922
rect 196 208894 3934 208908
rect 3962 208894 3967 208922
rect 297780 208418 298500 208516
rect 271777 208390 271782 208418
rect 271810 208404 298500 208418
rect 271810 208390 297836 208404
rect -480 201866 240 201964
rect -480 201852 6286 201866
rect 196 201838 6286 201852
rect 6314 201838 6319 201866
rect 297780 201810 298500 201908
rect 295465 201782 295470 201810
rect 295498 201796 298500 201810
rect 295498 201782 297836 201796
rect 297780 195202 298500 195300
rect 276761 195174 276766 195202
rect 276794 195188 298500 195202
rect 276794 195174 297836 195188
rect -480 194810 240 194908
rect -480 194796 6342 194810
rect 196 194782 6342 194796
rect 6370 194782 6375 194810
rect 297780 188594 298500 188692
rect 271833 188566 271838 188594
rect 271866 188580 298500 188594
rect 271866 188566 297836 188580
rect -480 187754 240 187852
rect -480 187740 4942 187754
rect 196 187726 4942 187740
rect 4970 187726 4975 187754
rect 297780 181986 298500 182084
rect 272729 181958 272734 181986
rect 272762 181972 298500 181986
rect 272762 181958 297836 181972
rect -480 180698 240 180796
rect -480 180684 2310 180698
rect 196 180670 2310 180684
rect 2338 180670 2343 180698
rect 297780 175378 298500 175476
rect 271889 175350 271894 175378
rect 271922 175364 298500 175378
rect 271922 175350 297836 175364
rect -480 173642 240 173740
rect -480 173628 3150 173642
rect 196 173614 3150 173628
rect 3178 173614 3183 173642
rect 297780 168770 298500 168868
rect 199481 168742 199486 168770
rect 199514 168742 205534 168770
rect 205562 168742 205567 168770
rect 271945 168742 271950 168770
rect 271978 168756 298500 168770
rect 271978 168742 297836 168756
rect 125561 168686 125566 168714
rect 125594 168686 135198 168714
rect 135226 168686 135231 168714
rect 198361 168686 198366 168714
rect 198394 168686 207046 168714
rect 207074 168686 207079 168714
rect 60265 168630 60270 168658
rect 60298 168630 69958 168658
rect 69986 168630 69991 168658
rect 114697 168630 114702 168658
rect 114730 168630 127134 168658
rect 127162 168630 127167 168658
rect 129929 168630 129934 168658
rect 129962 168630 143262 168658
rect 143290 168630 143295 168658
rect 191641 168630 191646 168658
rect 191674 168630 202062 168658
rect 202090 168630 202095 168658
rect 60937 168574 60942 168602
rect 60970 168574 71302 168602
rect 71330 168574 71335 168602
rect 116041 168574 116046 168602
rect 116074 168574 129822 168602
rect 129850 168574 129855 168602
rect 131609 168574 131614 168602
rect 131642 168574 145950 168602
rect 145978 168574 145983 168602
rect 180553 168574 180558 168602
rect 180586 168574 188846 168602
rect 188874 168574 188879 168602
rect 197241 168574 197246 168602
rect 197274 168574 207886 168602
rect 207914 168574 207919 168602
rect 63401 168518 63406 168546
rect 63434 168518 73990 168546
rect 74018 168518 74023 168546
rect 116713 168518 116718 168546
rect 116746 168518 131166 168546
rect 131194 168518 131199 168546
rect 132281 168518 132286 168546
rect 132314 168518 148638 168546
rect 148666 168518 148671 168546
rect 179881 168518 179886 168546
rect 179914 168518 188286 168546
rect 188314 168518 188319 168546
rect 193881 168518 193886 168546
rect 193914 168518 204750 168546
rect 204778 168518 204783 168546
rect 64409 168462 64414 168490
rect 64442 168462 75334 168490
rect 75362 168462 75367 168490
rect 117385 168462 117390 168490
rect 117418 168462 132510 168490
rect 132538 168462 132543 168490
rect 133961 168462 133966 168490
rect 133994 168462 151326 168490
rect 151354 168462 151359 168490
rect 179209 168462 179214 168490
rect 179242 168462 190526 168490
rect 190554 168462 190559 168490
rect 195001 168462 195006 168490
rect 195034 168462 206094 168490
rect 206122 168462 206127 168490
rect 22913 168406 22918 168434
rect 22946 168406 34062 168434
rect 34090 168406 34095 168434
rect 61609 168406 61614 168434
rect 61642 168406 72646 168434
rect 72674 168406 72679 168434
rect 118057 168406 118062 168434
rect 118090 168406 133854 168434
rect 133882 168406 133887 168434
rect 134969 168406 134974 168434
rect 135002 168406 154014 168434
rect 154042 168406 154047 168434
rect 175849 168406 175854 168434
rect 175882 168406 187726 168434
rect 187754 168406 187759 168434
rect 196121 168406 196126 168434
rect 196154 168406 207438 168434
rect 207466 168406 207471 168434
rect 254697 168406 254702 168434
rect 254730 168406 261198 168434
rect 261226 168406 261231 168434
rect 105289 168014 105294 168042
rect 105322 168014 109662 168042
rect 109690 168014 109695 168042
rect 239017 167958 239022 167986
rect 239050 167958 243950 167986
rect 243978 167958 243983 167986
rect 106633 167902 106638 167930
rect 106666 167902 112350 167930
rect 112378 167902 112383 167930
rect 240361 167902 240366 167930
rect 240394 167902 245294 167930
rect 245322 167902 245327 167930
rect 107305 167846 107310 167874
rect 107338 167846 113694 167874
rect 113722 167846 113727 167874
rect 241033 167846 241038 167874
rect 241066 167846 245966 167874
rect 245994 167846 245999 167874
rect 107977 167790 107982 167818
rect 108010 167790 115038 167818
rect 115066 167790 115071 167818
rect 50185 167734 50190 167762
rect 50218 167734 53830 167762
rect 53858 167734 53863 167762
rect 108649 167734 108654 167762
rect 108682 167734 116382 167762
rect 116410 167734 116415 167762
rect 236329 167734 236334 167762
rect 236362 167734 241262 167762
rect 241290 167734 241295 167762
rect 50857 167678 50862 167706
rect 50890 167678 55174 167706
rect 55202 167678 55207 167706
rect 109321 167678 109326 167706
rect 109354 167678 117726 167706
rect 117754 167678 117759 167706
rect 238345 167678 238350 167706
rect 238378 167678 243278 167706
rect 243306 167678 243311 167706
rect 109993 167622 109998 167650
rect 110026 167622 119070 167650
rect 119098 167622 119103 167650
rect 237001 167622 237006 167650
rect 237034 167622 241934 167650
rect 241962 167622 241967 167650
rect 52201 167566 52206 167594
rect 52234 167566 57862 167594
rect 57890 167566 57895 167594
rect 112009 167566 112014 167594
rect 112042 167566 121758 167594
rect 121786 167566 121791 167594
rect 174505 167566 174510 167594
rect 174538 167566 181006 167594
rect 181034 167566 181039 167594
rect 237673 167566 237678 167594
rect 237706 167566 242606 167594
rect 242634 167566 242639 167594
rect 103273 167342 103278 167370
rect 103306 167342 105630 167370
rect 105658 167342 105663 167370
rect 105961 167342 105966 167370
rect 105994 167342 111006 167370
rect 111034 167342 111039 167370
rect 102601 167286 102606 167314
rect 102634 167286 104286 167314
rect 104314 167286 104319 167314
rect 48169 167230 48174 167258
rect 48202 167230 49798 167258
rect 49826 167230 49831 167258
rect 181225 167230 181230 167258
rect 181258 167230 183806 167258
rect 183834 167230 183839 167258
rect 187945 167230 187950 167258
rect 187978 167230 189406 167258
rect 189434 167230 189439 167258
rect 47497 167174 47502 167202
rect 47530 167174 48454 167202
rect 48482 167174 48487 167202
rect 48841 167174 48846 167202
rect 48874 167174 51142 167202
rect 51170 167174 51175 167202
rect 51529 167174 51534 167202
rect 51562 167174 56518 167202
rect 56546 167174 56551 167202
rect 101929 167174 101934 167202
rect 101962 167174 102942 167202
rect 102970 167174 102975 167202
rect 181897 167174 181902 167202
rect 181930 167174 184366 167202
rect 184394 167174 184399 167202
rect 188617 167174 188622 167202
rect 188650 167174 189966 167202
rect 189994 167174 189999 167202
rect 239689 167174 239694 167202
rect 239722 167174 244622 167202
rect 244650 167174 244655 167202
rect 56905 167006 56910 167034
rect 56938 167006 63238 167034
rect 63266 167006 63271 167034
rect 57577 166950 57582 166978
rect 57610 166950 64582 166978
rect 64610 166950 64615 166978
rect 53545 166894 53550 166922
rect 53578 166894 60550 166922
rect 60578 166894 60583 166922
rect 58249 166838 58254 166866
rect 58282 166838 65926 166866
rect 65954 166838 65959 166866
rect 58921 166782 58926 166810
rect 58954 166782 67270 166810
rect 67298 166782 67303 166810
rect 26945 166726 26950 166754
rect 26978 166726 36078 166754
rect 36106 166726 36111 166754
rect 52873 166726 52878 166754
rect 52906 166726 59206 166754
rect 59234 166726 59239 166754
rect 59593 166726 59598 166754
rect 59626 166726 68614 166754
rect 68642 166726 68647 166754
rect 215105 166726 215110 166754
rect 215138 166726 223566 166754
rect 223594 166726 223599 166754
rect -480 166586 240 166684
rect -480 166572 3990 166586
rect 196 166558 3990 166572
rect 4018 166558 4023 166586
rect 235657 166278 235662 166306
rect 235690 166278 240590 166306
rect 240618 166278 240623 166306
rect 232969 166222 232974 166250
rect 233002 166222 237902 166250
rect 237930 166222 237935 166250
rect 234985 166166 234990 166194
rect 235018 166166 239918 166194
rect 239946 166166 239951 166194
rect 247977 165998 247982 166026
rect 248010 165998 254478 166026
rect 254506 165998 254511 166026
rect 232297 165942 232302 165970
rect 232330 165942 237230 165970
rect 237258 165942 237263 165970
rect 251337 165942 251342 165970
rect 251370 165942 257838 165970
rect 257866 165942 257871 165970
rect 175177 165886 175182 165914
rect 175210 165886 181566 165914
rect 181594 165886 181599 165914
rect 230281 165886 230286 165914
rect 230314 165886 235886 165914
rect 235914 165886 235919 165914
rect 248649 165886 248654 165914
rect 248682 165886 255150 165914
rect 255178 165886 255183 165914
rect 233641 165830 233646 165858
rect 233674 165830 238574 165858
rect 238602 165830 238607 165858
rect 234313 165774 234318 165802
rect 234346 165774 239246 165802
rect 239274 165774 239279 165802
rect 70961 165046 70966 165074
rect 70994 165046 80710 165074
rect 80738 165046 80743 165074
rect 253353 165046 253358 165074
rect 253386 165046 259854 165074
rect 259882 165046 259887 165074
rect 182121 164598 182126 164626
rect 182154 164598 182574 164626
rect 182602 164598 182607 164626
rect 182681 164598 182686 164626
rect 182714 164598 183246 164626
rect 183274 164598 183279 164626
rect 247305 164318 247310 164346
rect 247338 164318 253806 164346
rect 253834 164318 253839 164346
rect 249993 164262 249998 164290
rect 250026 164262 256494 164290
rect 256522 164262 256527 164290
rect 30977 164206 30982 164234
rect 31010 164206 38094 164234
rect 38122 164206 38127 164234
rect 246633 164206 246638 164234
rect 246666 164206 253134 164234
rect 253162 164206 253167 164234
rect 104617 163758 104622 163786
rect 104650 163758 108318 163786
rect 108346 163758 108351 163786
rect 116769 163758 116774 163786
rect 116802 163758 120414 163786
rect 120442 163758 120447 163786
rect 254025 163478 254030 163506
rect 254058 163478 260526 163506
rect 260554 163478 260559 163506
rect 103945 163422 103950 163450
rect 103978 163422 106974 163450
rect 107002 163422 107007 163450
rect 120073 163422 120078 163450
rect 120106 163422 137886 163450
rect 137914 163422 137919 163450
rect 249321 163422 249326 163450
rect 249354 163422 255822 163450
rect 255850 163422 255855 163450
rect 121417 163366 121422 163394
rect 121450 163366 140574 163394
rect 140602 163366 140607 163394
rect 250665 163366 250670 163394
rect 250698 163366 257166 163394
rect 257194 163366 257199 163394
rect 49513 162974 49518 163002
rect 49546 162974 52486 163002
rect 52514 162974 52519 163002
rect 130825 162862 130830 162890
rect 130858 162862 155358 162890
rect 155386 162862 155391 162890
rect 201161 162862 201166 162890
rect 201194 162862 213486 162890
rect 213514 162862 213519 162890
rect 131497 162806 131502 162834
rect 131530 162806 156702 162834
rect 156730 162806 156735 162834
rect 201721 162806 201726 162834
rect 201754 162806 214158 162834
rect 214186 162806 214191 162834
rect 132169 162750 132174 162778
rect 132202 162750 158046 162778
rect 158074 162750 158079 162778
rect 202281 162750 202286 162778
rect 202314 162750 214830 162778
rect 214858 162750 214863 162778
rect 132841 162694 132846 162722
rect 132874 162694 159390 162722
rect 159418 162694 159423 162722
rect 202841 162694 202846 162722
rect 202874 162694 215502 162722
rect 215530 162694 215535 162722
rect 127465 162638 127470 162666
rect 127498 162638 132286 162666
rect 132314 162638 132319 162666
rect 133513 162638 133518 162666
rect 133546 162638 160734 162666
rect 160762 162638 160767 162666
rect 197801 162638 197806 162666
rect 197834 162638 201166 162666
rect 201194 162638 201199 162666
rect 203401 162638 203406 162666
rect 203434 162638 216174 162666
rect 216202 162638 216207 162666
rect 128809 162582 128814 162610
rect 128842 162582 133966 162610
rect 133994 162582 133999 162610
rect 134185 162582 134190 162610
rect 134218 162582 162078 162610
rect 162106 162582 162111 162610
rect 208721 162582 208726 162610
rect 208754 162582 221550 162610
rect 221578 162582 221583 162610
rect 252681 162582 252686 162610
rect 252714 162582 259182 162610
rect 259210 162582 259215 162610
rect 32321 162526 32326 162554
rect 32354 162526 38766 162554
rect 38794 162526 38799 162554
rect 112681 162526 112686 162554
rect 112714 162526 123102 162554
rect 123130 162526 123135 162554
rect 126121 162526 126126 162554
rect 126154 162526 131614 162554
rect 131642 162526 131647 162554
rect 134857 162526 134862 162554
rect 134890 162526 163422 162554
rect 163450 162526 163455 162554
rect 198921 162526 198926 162554
rect 198954 162526 202454 162554
rect 202482 162526 202487 162554
rect 203961 162526 203966 162554
rect 203994 162526 216846 162554
rect 216874 162526 216879 162554
rect 252009 162526 252014 162554
rect 252042 162526 258510 162554
rect 258538 162526 258543 162554
rect 200041 162470 200046 162498
rect 200074 162470 203294 162498
rect 203322 162470 203327 162498
rect 200601 162414 200606 162442
rect 200634 162414 203518 162442
rect 203546 162414 203551 162442
rect 297780 162162 298500 162260
rect 41729 162134 41734 162162
rect 41762 162134 44142 162162
rect 44170 162134 44175 162162
rect 130153 162134 130158 162162
rect 130186 162134 134974 162162
rect 135002 162134 135007 162162
rect 272785 162134 272790 162162
rect 272818 162148 298500 162162
rect 272818 162134 297836 162148
rect 36353 162078 36358 162106
rect 36386 162078 40782 162106
rect 40810 162078 40815 162106
rect 44417 162078 44422 162106
rect 44450 162078 45486 162106
rect 45514 162078 45519 162106
rect 62281 162078 62286 162106
rect 62314 162078 63406 162106
rect 63434 162078 63439 162106
rect 86081 162078 86086 162106
rect 86114 162078 87822 162106
rect 87850 162078 87855 162106
rect 91849 162078 91854 162106
rect 91882 162078 93646 162106
rect 93674 162078 93679 162106
rect 118729 162078 118734 162106
rect 118762 162078 125566 162106
rect 125594 162078 125599 162106
rect 201161 162078 201166 162106
rect 201194 162078 209454 162106
rect 209482 162078 209487 162106
rect 62953 162022 62958 162050
rect 62986 162022 64414 162050
rect 64442 162022 64447 162050
rect 89833 162022 89838 162050
rect 89866 162022 93758 162050
rect 93786 162022 93791 162050
rect 119401 162022 119406 162050
rect 119434 162022 136542 162050
rect 136570 162022 136575 162050
rect 191081 162022 191086 162050
rect 191114 162022 201390 162050
rect 201418 162022 201423 162050
rect 202449 162022 202454 162050
rect 202482 162022 207046 162050
rect 207074 162022 207079 162050
rect 207153 162022 207158 162050
rect 207186 162022 210126 162050
rect 210154 162022 210159 162050
rect 65641 161966 65646 161994
rect 65674 161966 70966 161994
rect 70994 161966 70999 161994
rect 124105 161966 124110 161994
rect 124138 161966 141918 161994
rect 141946 161966 141951 161994
rect 192201 161966 192206 161994
rect 192234 161966 202734 161994
rect 202762 161966 202767 161994
rect 203289 161966 203294 161994
rect 203322 161966 212142 161994
rect 212170 161966 212175 161994
rect 63625 161910 63630 161938
rect 63658 161910 76678 161938
rect 76706 161910 76711 161938
rect 120745 161910 120750 161938
rect 120778 161910 139230 161938
rect 139258 161910 139263 161938
rect 192761 161910 192766 161938
rect 192794 161910 203406 161938
rect 203434 161910 203439 161938
rect 203513 161910 203518 161938
rect 203546 161910 212814 161938
rect 212842 161910 212847 161938
rect 29633 161854 29638 161882
rect 29666 161854 37422 161882
rect 37450 161854 37455 161882
rect 39041 161854 39046 161882
rect 39074 161854 42126 161882
rect 42154 161854 42159 161882
rect 64297 161854 64302 161882
rect 64330 161854 78022 161882
rect 78050 161854 78055 161882
rect 110665 161854 110670 161882
rect 110698 161854 116774 161882
rect 116802 161854 116807 161882
rect 125449 161854 125454 161882
rect 125482 161854 144606 161882
rect 144634 161854 144639 161882
rect 193321 161854 193326 161882
rect 193354 161854 204078 161882
rect 204106 161854 204111 161882
rect 28289 161798 28294 161826
rect 28322 161798 36750 161826
rect 36778 161798 36783 161826
rect 37697 161798 37702 161826
rect 37730 161798 41454 161826
rect 41482 161798 41487 161826
rect 64969 161798 64974 161826
rect 65002 161798 79366 161826
rect 79394 161798 79399 161826
rect 90505 161798 90510 161826
rect 90538 161798 95326 161826
rect 95354 161798 95359 161826
rect 113353 161798 113358 161826
rect 113386 161798 124446 161826
rect 124474 161798 124479 161826
rect 126793 161798 126798 161826
rect 126826 161798 147294 161826
rect 147322 161798 147327 161826
rect 194441 161798 194446 161826
rect 194474 161798 205422 161826
rect 205450 161798 205455 161826
rect 205529 161798 205534 161826
rect 205562 161798 211470 161826
rect 211498 161798 211503 161826
rect 25601 161742 25606 161770
rect 25634 161742 35406 161770
rect 35434 161742 35439 161770
rect 66313 161742 66318 161770
rect 66346 161742 82054 161770
rect 82082 161742 82087 161770
rect 93193 161742 93198 161770
rect 93226 161742 99638 161770
rect 99666 161742 99671 161770
rect 114025 161742 114030 161770
rect 114058 161742 125790 161770
rect 125818 161742 125823 161770
rect 128137 161742 128142 161770
rect 128170 161742 149982 161770
rect 150010 161742 150015 161770
rect 195561 161742 195566 161770
rect 195594 161742 206766 161770
rect 206794 161742 206799 161770
rect 207041 161742 207046 161770
rect 207074 161742 210798 161770
rect 210826 161742 210831 161770
rect 216281 161742 216286 161770
rect 216314 161742 222222 161770
rect 222250 161742 222255 161770
rect 24257 161686 24262 161714
rect 24290 161686 34734 161714
rect 34762 161686 34767 161714
rect 35009 161686 35014 161714
rect 35042 161686 40110 161714
rect 40138 161686 40143 161714
rect 56233 161686 56238 161714
rect 56266 161686 61894 161714
rect 61922 161686 61927 161714
rect 66985 161686 66990 161714
rect 67018 161686 83398 161714
rect 83426 161686 83431 161714
rect 91177 161686 91182 161714
rect 91210 161686 99526 161714
rect 99554 161686 99559 161714
rect 115369 161686 115374 161714
rect 115402 161686 128478 161714
rect 128506 161686 128511 161714
rect 129481 161686 129486 161714
rect 129514 161686 152670 161714
rect 152698 161686 152703 161714
rect 196681 161686 196686 161714
rect 196714 161686 208110 161714
rect 208138 161686 208143 161714
rect 216393 161686 216398 161714
rect 216426 161686 222894 161714
rect 222922 161686 222927 161714
rect 230953 161686 230958 161714
rect 230986 161686 236558 161714
rect 236586 161686 236591 161714
rect 124777 161630 124782 161658
rect 124810 161630 129934 161658
rect 129962 161630 129967 161658
rect 86921 161350 86926 161378
rect 86954 161350 89166 161378
rect 89194 161350 89199 161378
rect 33665 161294 33670 161322
rect 33698 161294 39438 161322
rect 39466 161294 39471 161322
rect 40385 161294 40390 161322
rect 40418 161294 42798 161322
rect 42826 161294 42831 161322
rect 43073 161294 43078 161322
rect 43106 161294 44814 161322
rect 44842 161294 44847 161322
rect 87033 161294 87038 161322
rect 87066 161294 88494 161322
rect 88522 161294 88527 161322
rect 92521 161294 92526 161322
rect 92554 161294 95438 161322
rect 95466 161294 95471 161322
rect 207881 161294 207886 161322
rect 207914 161294 208782 161322
rect 208810 161294 208815 161322
rect 216505 161294 216510 161322
rect 216538 161294 220878 161322
rect 220906 161294 220911 161322
rect 224233 161294 224238 161322
rect 224266 161294 224686 161322
rect 224714 161294 224719 161322
rect 224905 161294 224910 161322
rect 224938 161294 227206 161322
rect 227234 161294 227239 161322
rect -480 159530 240 159628
rect -480 159516 6398 159530
rect 196 159502 6398 159516
rect 6426 159502 6431 159530
rect 269705 159334 269710 159362
rect 269738 159334 269743 159362
rect 269710 159012 269738 159334
rect 269948 158550 273406 158578
rect 273434 158550 273439 158578
rect 269948 158102 292334 158130
rect 292362 158102 292367 158130
rect 20393 157766 20398 157794
rect 20426 157766 30044 157794
rect 269948 157654 275926 157682
rect 275954 157654 275959 157682
rect 16529 157206 16534 157234
rect 16562 157206 30044 157234
rect 269948 157206 271726 157234
rect 271754 157206 271759 157234
rect 269948 156758 295246 156786
rect 295274 156758 295279 156786
rect 5497 156646 5502 156674
rect 5530 156646 30044 156674
rect 269948 156310 275086 156338
rect 275114 156310 275119 156338
rect 3761 156086 3766 156114
rect 3794 156086 30044 156114
rect 269948 155862 278446 155890
rect 278474 155862 278479 155890
rect 297780 155554 298500 155652
rect 2081 155526 2086 155554
rect 2114 155526 30044 155554
rect 271721 155526 271726 155554
rect 271754 155540 298500 155554
rect 271754 155526 297836 155540
rect 269948 155414 295302 155442
rect 295330 155414 295335 155442
rect 5441 154966 5446 154994
rect 5474 154966 30044 154994
rect 269948 154966 272566 154994
rect 272594 154966 272599 154994
rect 269948 154518 272622 154546
rect 272650 154518 272655 154546
rect 3089 154406 3094 154434
rect 3122 154406 30044 154434
rect 269948 154070 295358 154098
rect 295386 154070 295391 154098
rect 2137 153846 2142 153874
rect 2170 153846 30044 153874
rect 269948 153622 273406 153650
rect 273434 153622 273439 153650
rect 5497 153286 5502 153314
rect 5530 153286 30044 153314
rect 269948 153174 277606 153202
rect 277634 153174 277639 153202
rect 3817 152726 3822 152754
rect 3850 152726 30044 152754
rect 269948 152726 295414 152754
rect 295442 152726 295447 152754
rect -480 152474 240 152572
rect -480 152460 2086 152474
rect 196 152446 2086 152460
rect 2114 152446 2119 152474
rect 269948 152278 272678 152306
rect 272706 152278 272711 152306
rect 2193 152166 2198 152194
rect 2226 152166 30044 152194
rect 269948 151830 271782 151858
rect 271810 151830 271815 151858
rect 5553 151606 5558 151634
rect 5586 151606 30044 151634
rect 269948 151382 295470 151410
rect 295498 151382 295503 151410
rect 3873 151046 3878 151074
rect 3906 151046 30044 151074
rect 269948 150934 276766 150962
rect 276794 150934 276799 150962
rect 2249 150486 2254 150514
rect 2282 150486 30044 150514
rect 269948 150486 271838 150514
rect 271866 150486 271871 150514
rect 269948 150038 272734 150066
rect 272762 150038 272767 150066
rect 5609 149926 5614 149954
rect 5642 149926 30044 149954
rect 269948 149590 271894 149618
rect 271922 149590 271927 149618
rect 3929 149366 3934 149394
rect 3962 149366 30044 149394
rect 269948 149142 271950 149170
rect 271978 149142 271983 149170
rect 297780 148932 298500 149044
rect 6281 148806 6286 148834
rect 6314 148806 30044 148834
rect 269948 148694 272790 148722
rect 272818 148694 272823 148722
rect 6337 148246 6342 148274
rect 6370 148246 30044 148274
rect 269948 148246 271726 148274
rect 271754 148246 271759 148274
rect 4937 147686 4942 147714
rect 4970 147686 30044 147714
rect 269948 147350 271894 147378
rect 271922 147350 271927 147378
rect 2305 147126 2310 147154
rect 2338 147126 30044 147154
rect 269948 146902 271782 146930
rect 271810 146902 271815 146930
rect 3145 146566 3150 146594
rect 3178 146566 30044 146594
rect 3985 146006 3990 146034
rect 4018 146006 30044 146034
rect 269948 146006 276990 146034
rect 277018 146006 277023 146034
rect 269948 145558 271726 145586
rect 271754 145558 271759 145586
rect -480 145418 240 145516
rect 6393 145446 6398 145474
rect 6426 145446 30044 145474
rect -480 145404 2478 145418
rect 196 145390 2478 145404
rect 2506 145390 2511 145418
rect 2081 144886 2086 144914
rect 2114 144886 30044 144914
rect 269948 144662 276934 144690
rect 276962 144662 276967 144690
rect 2473 144326 2478 144354
rect 2506 144326 30044 144354
rect 269948 144214 271838 144242
rect 271866 144214 271871 144242
rect 2081 143766 2086 143794
rect 2114 143766 30044 143794
rect 269948 143318 276878 143346
rect 276906 143318 276911 143346
rect 28233 143206 28238 143234
rect 28266 143206 30044 143234
rect 269948 142870 271950 142898
rect 271978 142870 271983 142898
rect 28177 142646 28182 142674
rect 28210 142646 30044 142674
rect 297780 142338 298500 142436
rect 271889 142310 271894 142338
rect 271922 142324 298500 142338
rect 271922 142310 297836 142324
rect 2361 142086 2366 142114
rect 2394 142086 30044 142114
rect 269948 141974 276150 142002
rect 276178 141974 276183 142002
rect 28121 141526 28126 141554
rect 28154 141526 30044 141554
rect 269948 141526 276822 141554
rect 276850 141526 276855 141554
rect 3145 140966 3150 140994
rect 3178 140966 30044 140994
rect 269948 140630 276038 140658
rect 276066 140630 276071 140658
rect 6281 140406 6286 140434
rect 6314 140406 30044 140434
rect 269948 140182 276766 140210
rect 276794 140182 276799 140210
rect 3985 139846 3990 139874
rect 4018 139846 30044 139874
rect 3929 139286 3934 139314
rect 3962 139286 30044 139314
rect 269948 139286 276094 139314
rect 276122 139286 276127 139314
rect 269948 138838 275982 138866
rect 276010 138838 276015 138866
rect 7121 138726 7126 138754
rect 7154 138726 30044 138754
rect 196 138460 2086 138474
rect -480 138446 2086 138460
rect 2114 138446 2119 138474
rect -480 138348 240 138446
rect 2305 138166 2310 138194
rect 2338 138166 30044 138194
rect 269948 137942 275926 137970
rect 275954 137942 275959 137970
rect 3873 137606 3878 137634
rect 3906 137606 30044 137634
rect 269948 137494 277606 137522
rect 277634 137494 277639 137522
rect 2249 137046 2254 137074
rect 2282 137046 30044 137074
rect 269948 137046 277718 137074
rect 277746 137046 277751 137074
rect 269948 136598 277830 136626
rect 277858 136598 277863 136626
rect 2193 136486 2198 136514
rect 2226 136486 30044 136514
rect 269948 136150 277942 136178
rect 277970 136150 277975 136178
rect 3089 135926 3094 135954
rect 3122 135926 30044 135954
rect 297780 135730 298500 135828
rect 269934 135674 269962 135716
rect 271777 135702 271782 135730
rect 271810 135716 298500 135730
rect 271810 135702 297836 135716
rect 269934 135646 275422 135674
rect 275450 135646 275455 135674
rect 3817 135366 3822 135394
rect 3850 135366 30044 135394
rect 269948 135254 272118 135282
rect 272146 135254 272151 135282
rect 5441 134806 5446 134834
rect 5474 134806 30044 134834
rect 269948 134806 278166 134834
rect 278194 134806 278199 134834
rect 269948 134358 276430 134386
rect 276458 134358 276463 134386
rect 3761 134246 3766 134274
rect 3794 134246 30044 134274
rect 269948 133910 276374 133938
rect 276402 133910 276407 133938
rect 2137 133686 2142 133714
rect 2170 133686 30044 133714
rect 269948 133462 278222 133490
rect 278250 133462 278255 133490
rect 2081 133126 2086 133154
rect 2114 133126 30044 133154
rect 269948 133014 275590 133042
rect 275618 133014 275623 133042
rect 21401 132566 21406 132594
rect 21434 132566 30044 132594
rect 269948 132566 275646 132594
rect 275674 132566 275679 132594
rect 269948 132118 278054 132146
rect 278082 132118 278087 132146
rect 19273 132006 19278 132034
rect 19306 132006 30044 132034
rect 269948 131670 277214 131698
rect 277242 131670 277247 131698
rect -480 131306 240 131404
rect -480 131292 28238 131306
rect 196 131278 28238 131292
rect 28266 131278 28271 131306
rect 269948 131222 278110 131250
rect 278138 131222 278143 131250
rect 269948 130774 278278 130802
rect 278306 130774 278311 130802
rect 97561 129318 97566 129346
rect 97594 129318 102886 129346
rect 102914 129318 102919 129346
rect 124665 129318 124670 129346
rect 124698 129318 132510 129346
rect 132538 129318 132543 129346
rect 236665 129318 236670 129346
rect 236698 129318 245014 129346
rect 245042 129318 245047 129346
rect 95545 129262 95550 129290
rect 95578 129262 102438 129290
rect 102466 129262 102471 129290
rect 118617 129262 118622 129290
rect 118650 129262 126462 129290
rect 126490 129262 126495 129290
rect 126681 129262 126686 129290
rect 126714 129262 134526 129290
rect 134554 129262 134559 129290
rect 233305 129262 233310 129290
rect 233338 129262 242718 129290
rect 242746 129262 242751 129290
rect 61945 129206 61950 129234
rect 61978 129206 66990 129234
rect 67018 129206 67023 129234
rect 91513 129206 91518 129234
rect 91546 129206 99134 129234
rect 99162 129206 99167 129234
rect 100921 129206 100926 129234
rect 100954 129206 107870 129234
rect 107898 129206 107903 129234
rect 121305 129206 121310 129234
rect 121338 129206 129150 129234
rect 129178 129206 129183 129234
rect 223225 129206 223230 129234
rect 223258 129206 230958 129234
rect 230986 129206 230991 129234
rect 233977 129206 233982 129234
rect 234010 129206 243558 129234
rect 243586 129206 243591 129234
rect 66761 129150 66766 129178
rect 66794 129150 76062 129178
rect 76090 129150 76095 129178
rect 96889 129150 96894 129178
rect 96922 129150 106526 129178
rect 106554 129150 106559 129178
rect 119289 129150 119294 129178
rect 119322 129150 127134 129178
rect 127162 129150 127167 129178
rect 224569 129150 224574 129178
rect 224602 129150 232246 129178
rect 232274 129150 232279 129178
rect 241369 129150 241374 129178
rect 241402 129150 251566 129178
rect 251594 129150 251599 129178
rect 55897 129094 55902 129122
rect 55930 129094 68446 129122
rect 68474 129094 68479 129122
rect 98233 129094 98238 129122
rect 98266 129094 110054 129122
rect 110082 129094 110087 129122
rect 121977 129094 121982 129122
rect 122010 129094 129822 129122
rect 129850 129094 129855 129122
rect 172097 129094 172102 129122
rect 172130 129094 178878 129122
rect 178906 129094 178911 129122
rect 179937 129094 179942 129122
rect 179970 129094 183582 129122
rect 183610 129094 183615 129122
rect 203737 129094 203742 129122
rect 203770 129094 213542 129122
rect 213570 129094 213575 129122
rect 222553 129094 222558 129122
rect 222586 129094 231798 129122
rect 231826 129094 231831 129122
rect 234649 129094 234654 129122
rect 234682 129094 258342 129122
rect 258370 129094 258375 129122
rect 297780 129108 298500 129220
rect 33945 129038 33950 129066
rect 33978 129038 41790 129066
rect 41818 129038 41823 129066
rect 53881 129038 53886 129066
rect 53914 129038 66878 129066
rect 66906 129038 66911 129066
rect 70121 129038 70126 129066
rect 70154 129038 76734 129066
rect 76762 129038 76767 129066
rect 94201 129038 94206 129066
rect 94234 129038 109046 129066
rect 109074 129038 109079 129066
rect 114585 129038 114590 129066
rect 114618 129038 121086 129066
rect 121114 129038 121119 129066
rect 126009 129038 126014 129066
rect 126042 129038 133854 129066
rect 133882 129038 133887 129066
rect 170977 129038 170982 129066
rect 171010 129038 178206 129066
rect 178234 129038 178239 129066
rect 178817 129038 178822 129066
rect 178850 129038 182910 129066
rect 182938 129038 182943 129066
rect 195673 129038 195678 129066
rect 195706 129038 200102 129066
rect 200130 129038 200135 129066
rect 210457 129038 210462 129066
rect 210490 129038 224742 129066
rect 224770 129038 224775 129066
rect 235993 129038 235998 129066
rect 236026 129038 260582 129066
rect 260610 129038 260615 129066
rect 16809 128982 16814 129010
rect 16842 128982 35070 129010
rect 35098 128982 35103 129010
rect 37361 128982 37366 129010
rect 37394 128982 72030 129010
rect 72058 128982 72063 129010
rect 90169 128982 90174 129010
rect 90202 128982 106806 129010
rect 106834 128982 106839 129010
rect 115257 128982 115262 129010
rect 115290 128982 123102 129010
rect 123130 128982 123135 129010
rect 127353 128982 127358 129010
rect 127386 128982 135198 129010
rect 135226 128982 135231 129010
rect 137993 128982 137998 129010
rect 138026 128982 144606 129010
rect 144634 128982 144639 129010
rect 148633 128982 148638 129010
rect 148666 128982 155134 129010
rect 155162 128982 155167 129010
rect 169857 128982 169862 129010
rect 169890 128982 177534 129010
rect 177562 128982 177567 129010
rect 196345 128982 196350 129010
rect 196378 128982 201222 129010
rect 201250 128982 201255 129010
rect 211801 128982 211806 129010
rect 211834 128982 226982 129010
rect 227010 128982 227015 129010
rect 232633 128982 232638 129010
rect 232666 128982 239414 129010
rect 239442 128982 239447 129010
rect 240025 128982 240030 129010
rect 240058 128982 265398 129010
rect 265426 128982 265431 129010
rect 34841 128926 34846 128954
rect 34874 128926 70686 128954
rect 70714 128926 70719 128954
rect 86137 128926 86142 128954
rect 86170 128926 108150 128954
rect 108178 128926 108183 128954
rect 115929 128926 115934 128954
rect 115962 128926 123774 128954
rect 123802 128926 123807 128954
rect 132281 128926 132286 128954
rect 132314 128926 143262 128954
rect 143290 128926 143295 128954
rect 149977 128926 149982 128954
rect 150010 128926 159166 128954
rect 159194 128926 159199 128954
rect 163137 128926 163142 128954
rect 163170 128926 173502 128954
rect 173530 128926 173535 128954
rect 174337 128926 174342 128954
rect 174370 128926 180222 128954
rect 180250 128926 180255 128954
rect 182177 128926 182182 128954
rect 182210 128926 184926 128954
rect 184954 128926 184959 128954
rect 197017 128926 197022 128954
rect 197050 128926 202342 128954
rect 202370 128926 202375 128954
rect 204409 128926 204414 128954
rect 204442 128926 214662 128954
rect 214690 128926 214695 128954
rect 217849 128926 217854 128954
rect 217882 128926 233814 128954
rect 233842 128926 233847 128954
rect 237337 128926 237342 128954
rect 237370 128926 262822 128954
rect 262850 128926 262855 128954
rect 47833 128870 47838 128898
rect 47866 128870 48286 128898
rect 48314 128870 48319 128898
rect 49177 128870 49182 128898
rect 49210 128870 49966 128898
rect 49994 128870 49999 128898
rect 75833 128870 75838 128898
rect 75866 128870 77406 128898
rect 77434 128870 77439 128898
rect 112569 128870 112574 128898
rect 112602 128870 115038 128898
rect 115066 128870 115071 128898
rect 117721 128870 117726 128898
rect 117754 128870 118846 128898
rect 118874 128870 118879 128898
rect 120633 128870 120638 128898
rect 120666 128870 128478 128898
rect 128506 128870 128511 128898
rect 181057 128870 181062 128898
rect 181090 128870 184254 128898
rect 184282 128870 184287 128898
rect 184417 128870 184422 128898
rect 184450 128870 186270 128898
rect 186298 128870 186303 128898
rect 190297 128870 190302 128898
rect 190330 128870 191142 128898
rect 191170 128870 191175 128898
rect 118393 128814 118398 128842
rect 118426 128814 119070 128842
rect 119098 128814 119103 128842
rect 183297 128814 183302 128842
rect 183330 128814 185598 128842
rect 185626 128814 185631 128842
rect 190969 128814 190974 128842
rect 191002 128814 192262 128842
rect 192290 128814 192295 128842
rect 112345 128646 112350 128674
rect 112378 128646 116886 128674
rect 116914 128646 116919 128674
rect 113241 128590 113246 128618
rect 113274 128590 117054 128618
rect 117082 128590 117087 128618
rect 51193 128534 51198 128562
rect 51226 128534 51646 128562
rect 51674 128534 51679 128562
rect 120521 128534 120526 128562
rect 120554 128534 122430 128562
rect 122458 128534 122463 128562
rect 177697 128534 177702 128562
rect 177730 128534 182238 128562
rect 182266 128534 182271 128562
rect 185537 128534 185542 128562
rect 185570 128534 186942 128562
rect 186970 128534 186975 128562
rect 223897 128534 223902 128562
rect 223930 128534 228494 128562
rect 228522 128534 228527 128562
rect 106801 128478 106806 128506
rect 106834 128478 109494 128506
rect 109522 128478 109527 128506
rect 239386 128478 250502 128506
rect 250530 128478 250535 128506
rect 98905 128366 98910 128394
rect 98938 128366 107198 128394
rect 107226 128366 107231 128394
rect 239386 128338 239414 128478
rect 106297 128310 106302 128338
rect 106330 128310 115038 128338
rect 115066 128310 115071 128338
rect 229945 128310 229950 128338
rect 229978 128310 239414 128338
rect 247870 128422 251622 128450
rect 251650 128422 251655 128450
rect 247870 128282 247898 128422
rect 101593 128254 101598 128282
rect 101626 128254 113470 128282
rect 113498 128254 113503 128282
rect 230617 128254 230622 128282
rect 230650 128254 247898 128282
rect 247926 128310 248290 128338
rect 247926 128226 247954 128310
rect 248262 128282 248290 128310
rect 248262 128254 248654 128282
rect 251561 128254 251566 128282
rect 251594 128254 269542 128282
rect 269570 128254 269575 128282
rect 99577 128198 99582 128226
rect 99610 128198 112798 128226
rect 112826 128198 112831 128226
rect 231289 128198 231294 128226
rect 231322 128198 247954 128226
rect 248626 128226 248654 128254
rect 248626 128198 252770 128226
rect 252742 128170 252770 128198
rect 93529 128142 93534 128170
rect 93562 128142 110782 128170
rect 110810 128142 110815 128170
rect 111673 128142 111678 128170
rect 111706 128142 116830 128170
rect 116858 128142 116863 128170
rect 197689 128142 197694 128170
rect 197722 128142 203462 128170
rect 203490 128142 203495 128170
rect 231961 128142 231966 128170
rect 231994 128142 251370 128170
rect 252737 128142 252742 128170
rect 252770 128142 252775 128170
rect 89497 128086 89502 128114
rect 89530 128086 109438 128114
rect 109466 128086 109471 128114
rect 116601 128086 116606 128114
rect 116634 128086 124446 128114
rect 124474 128086 124479 128114
rect 175457 128086 175462 128114
rect 175490 128086 180894 128114
rect 180922 128086 180927 128114
rect 198361 128086 198366 128114
rect 198394 128086 204582 128114
rect 204610 128086 204615 128114
rect 212473 128086 212478 128114
rect 212506 128086 228102 128114
rect 228130 128086 228135 128114
rect 235321 128086 235326 128114
rect 235354 128086 248654 128114
rect 248626 128002 248654 128086
rect 251342 128058 251370 128142
rect 254506 128086 259462 128114
rect 259490 128086 259495 128114
rect 251342 128030 253862 128058
rect 253890 128030 253895 128058
rect 254506 128002 254534 128086
rect 248626 127974 254534 128002
rect 102881 127638 102886 127666
rect 102914 127638 112126 127666
rect 112154 127638 112159 127666
rect 242713 127638 242718 127666
rect 242746 127638 256102 127666
rect 256130 127638 256135 127666
rect 102433 127582 102438 127610
rect 102466 127582 111454 127610
rect 111482 127582 111487 127610
rect 239409 127582 239414 127610
rect 239442 127582 254982 127610
rect 255010 127582 255015 127610
rect 99129 127526 99134 127554
rect 99162 127526 110110 127554
rect 110138 127526 110143 127554
rect 203065 127526 203070 127554
rect 203098 127526 212422 127554
rect 212450 127526 212455 127554
rect 225241 127526 225246 127554
rect 225274 127526 242662 127554
rect 242690 127526 242695 127554
rect 243553 127526 243558 127554
rect 243586 127526 257222 127554
rect 257250 127526 257255 127554
rect 92857 127470 92862 127498
rect 92890 127470 105182 127498
rect 105210 127470 105215 127498
rect 109657 127470 109662 127498
rect 109690 127470 116158 127498
rect 116186 127470 116191 127498
rect 207769 127470 207774 127498
rect 207802 127470 220262 127498
rect 220290 127470 220295 127498
rect 226585 127470 226590 127498
rect 226618 127470 244902 127498
rect 244930 127470 244935 127498
rect 245009 127470 245014 127498
rect 245042 127470 261702 127498
rect 261730 127470 261735 127498
rect 88825 127414 88830 127442
rect 88858 127414 103838 127442
rect 103866 127414 103871 127442
rect 108313 127414 108318 127442
rect 108346 127414 115542 127442
rect 115570 127414 115575 127442
rect 208441 127414 208446 127442
rect 208474 127414 221382 127442
rect 221410 127414 221415 127442
rect 227257 127414 227262 127442
rect 227290 127414 246022 127442
rect 246050 127414 246055 127442
rect 86809 127358 86814 127386
rect 86842 127358 103166 127386
rect 103194 127358 103199 127386
rect 107641 127358 107646 127386
rect 107674 127358 115486 127386
rect 115514 127358 115519 127386
rect 209113 127358 209118 127386
rect 209146 127358 222502 127386
rect 222530 127358 222535 127386
rect 227929 127358 227934 127386
rect 227962 127358 247142 127386
rect 247170 127358 247175 127386
rect 84793 127302 84798 127330
rect 84826 127302 102494 127330
rect 102522 127302 102527 127330
rect 105625 127302 105630 127330
rect 105658 127302 114814 127330
rect 114842 127302 114847 127330
rect 199705 127302 199710 127330
rect 199738 127302 206822 127330
rect 206850 127302 206855 127330
rect 209785 127302 209790 127330
rect 209818 127302 223622 127330
rect 223650 127302 223655 127330
rect 228601 127302 228606 127330
rect 228634 127302 248262 127330
rect 248290 127302 248295 127330
rect 82777 127246 82782 127274
rect 82810 127246 102046 127274
rect 102074 127246 102079 127274
rect 102265 127246 102270 127274
rect 102298 127246 113694 127274
rect 113722 127246 113727 127274
rect 201721 127246 201726 127274
rect 201754 127246 210182 127274
rect 210210 127246 210215 127274
rect 211129 127246 211134 127274
rect 211162 127246 225862 127274
rect 225890 127246 225895 127274
rect 229273 127246 229278 127274
rect 229306 127246 249382 127274
rect 249410 127246 249415 127274
rect 102937 127190 102942 127218
rect 102970 127190 108542 127218
rect 108570 127190 108575 127218
rect 120185 126910 120190 126938
rect 120218 126910 121758 126938
rect 121786 126910 121791 126938
rect 104953 126854 104958 126882
rect 104986 126854 109214 126882
rect 109242 126854 109247 126882
rect 111897 126854 111902 126882
rect 111930 126854 113022 126882
rect 113050 126854 113055 126882
rect 119737 126854 119742 126882
rect 119770 126854 120414 126882
rect 120442 126854 120447 126882
rect 186657 126854 186662 126882
rect 186690 126854 187614 126882
rect 187642 126854 187647 126882
rect 100249 126798 100254 126826
rect 100282 126798 112854 126826
rect 112882 126798 112887 126826
rect 113745 126798 113750 126826
rect 113778 126798 117502 126826
rect 117530 126798 117535 126826
rect 176577 126798 176582 126826
rect 176610 126798 181566 126826
rect 181594 126798 181599 126826
rect 191641 126798 191646 126826
rect 191674 126798 193382 126826
rect 193410 126798 193415 126826
rect 207097 126798 207102 126826
rect 207130 126798 219142 126826
rect 219170 126798 219175 126826
rect 225913 126798 225918 126826
rect 225946 126798 243782 126826
rect 243810 126798 243815 126826
rect 90841 126742 90846 126770
rect 90874 126742 104510 126770
rect 104538 126742 104543 126770
rect 108985 126742 108990 126770
rect 109018 126742 110558 126770
rect 110586 126742 110591 126770
rect 195001 126742 195006 126770
rect 195034 126742 198982 126770
rect 199010 126742 199015 126770
rect 213145 126742 213150 126770
rect 213178 126742 229222 126770
rect 229250 126742 229255 126770
rect 238009 126742 238014 126770
rect 238042 126742 263942 126770
rect 263970 126742 263975 126770
rect 96217 126686 96222 126714
rect 96250 126686 107086 126714
rect 107114 126686 107119 126714
rect 119961 126686 119966 126714
rect 119994 126686 127806 126714
rect 127834 126686 127839 126714
rect 199033 126686 199038 126714
rect 199066 126686 205702 126714
rect 205730 126686 205735 126714
rect 213817 126686 213822 126714
rect 213850 126686 230342 126714
rect 230370 126686 230375 126714
rect 238681 126686 238686 126714
rect 238714 126686 265062 126714
rect 265090 126686 265095 126714
rect 92185 126630 92190 126658
rect 92218 126630 110334 126658
rect 110362 126630 110367 126658
rect 115705 126630 115710 126658
rect 115738 126630 118174 126658
rect 118202 126630 118207 126658
rect 122649 126630 122654 126658
rect 122682 126630 130494 126658
rect 130522 126630 130527 126658
rect 200377 126630 200382 126658
rect 200410 126630 207942 126658
rect 207970 126630 207975 126658
rect 214489 126630 214494 126658
rect 214522 126630 231462 126658
rect 231490 126630 231495 126658
rect 231793 126630 231798 126658
rect 231826 126630 238182 126658
rect 238210 126630 238215 126658
rect 239353 126630 239358 126658
rect 239386 126630 266182 126658
rect 266210 126630 266215 126658
rect 83449 126574 83454 126602
rect 83482 126574 102270 126602
rect 102298 126574 102303 126602
rect 103609 126574 103614 126602
rect 103642 126574 114142 126602
rect 114170 126574 114175 126602
rect 114361 126574 114366 126602
rect 114394 126574 117726 126602
rect 117754 126574 117759 126602
rect 117945 126574 117950 126602
rect 117978 126574 125790 126602
rect 125818 126574 125823 126602
rect 127666 126574 131166 126602
rect 131194 126574 131199 126602
rect 173217 126574 173222 126602
rect 173250 126574 179550 126602
rect 179578 126574 179583 126602
rect 201049 126574 201054 126602
rect 201082 126574 209062 126602
rect 209090 126574 209095 126602
rect 215161 126574 215166 126602
rect 215194 126574 232582 126602
rect 232610 126574 232615 126602
rect 240697 126574 240702 126602
rect 240730 126574 268422 126602
rect 268450 126574 268455 126602
rect 127666 126546 127694 126574
rect 88153 126518 88158 126546
rect 88186 126518 108990 126546
rect 109018 126518 109023 126546
rect 116377 126518 116382 126546
rect 116410 126518 118398 126546
rect 118426 126518 118431 126546
rect 123321 126518 123326 126546
rect 123354 126518 127694 126546
rect 168737 126518 168742 126546
rect 168770 126518 176862 126546
rect 176890 126518 176895 126546
rect 202393 126518 202398 126546
rect 202426 126518 211302 126546
rect 211330 126518 211335 126546
rect 215833 126518 215838 126546
rect 215866 126518 233702 126546
rect 233730 126518 233735 126546
rect 242041 126518 242046 126546
rect 242074 126518 270662 126546
rect 270690 126518 270695 126546
rect 87481 126462 87486 126490
rect 87514 126462 108766 126490
rect 108794 126462 108799 126490
rect 109041 126462 109046 126490
rect 109074 126462 111006 126490
rect 111034 126462 111039 126490
rect 113913 126462 113918 126490
rect 113946 126462 119014 126490
rect 119042 126462 119047 126490
rect 123993 126462 123998 126490
rect 124026 126462 131838 126490
rect 131866 126462 131871 126490
rect 167617 126462 167622 126490
rect 167650 126462 176190 126490
rect 176218 126462 176223 126490
rect 205081 126462 205086 126490
rect 205114 126462 215782 126490
rect 215810 126462 215815 126490
rect 216505 126462 216510 126490
rect 216538 126462 234822 126490
rect 234850 126462 234855 126490
rect 242601 126462 242606 126490
rect 242634 126462 271782 126490
rect 271810 126462 271815 126490
rect 85465 126406 85470 126434
rect 85498 126406 108094 126434
rect 108122 126406 108127 126434
rect 110385 126406 110390 126434
rect 110418 126406 116382 126434
rect 116410 126406 116415 126434
rect 117273 126406 117278 126434
rect 117306 126406 125118 126434
rect 125146 126406 125151 126434
rect 125337 126406 125342 126434
rect 125370 126406 133182 126434
rect 133210 126406 133215 126434
rect 166497 126406 166502 126434
rect 166530 126406 175518 126434
rect 175546 126406 175551 126434
rect 192313 126406 192318 126434
rect 192346 126406 194502 126434
rect 194530 126406 194535 126434
rect 205753 126406 205758 126434
rect 205786 126406 216902 126434
rect 216930 126406 216935 126434
rect 217177 126406 217182 126434
rect 217210 126406 235942 126434
rect 235970 126406 235975 126434
rect 243385 126406 243390 126434
rect 243418 126406 272902 126434
rect 272930 126406 272935 126434
rect 94873 126350 94878 126378
rect 94906 126350 105854 126378
rect 105882 126350 105887 126378
rect 107081 126350 107086 126378
rect 107114 126350 111678 126378
rect 111706 126350 111711 126378
rect 206425 126350 206430 126378
rect 206458 126350 218022 126378
rect 218050 126350 218055 126378
rect 228489 126350 228494 126378
rect 228522 126350 240422 126378
rect 240450 126350 240455 126378
rect 104281 126294 104286 126322
rect 104314 126294 114366 126322
rect 114394 126294 114399 126322
rect 232241 126294 232246 126322
rect 232274 126294 241542 126322
rect 241570 126294 241575 126322
rect 192985 126238 192990 126266
rect 193018 126238 195622 126266
rect 195650 126238 195655 126266
rect 230953 126238 230958 126266
rect 230986 126238 239302 126266
rect 239330 126238 239335 126266
rect 193657 126182 193662 126210
rect 193690 126182 196742 126210
rect 196770 126182 196775 126210
rect 233809 126182 233814 126210
rect 233842 126182 237062 126210
rect 237090 126182 237095 126210
rect 265393 126182 265398 126210
rect 265426 126182 267302 126210
rect 267330 126182 267335 126210
rect 106969 126126 106974 126154
rect 107002 126126 109886 126154
rect 109914 126126 109919 126154
rect 110049 126126 110054 126154
rect 110082 126126 112350 126154
rect 112378 126126 112383 126154
rect 194329 126126 194334 126154
rect 194362 126126 197862 126154
rect 197890 126126 197895 126154
rect 271945 125678 271950 125706
rect 271978 125678 295246 125706
rect 295274 125678 295279 125706
rect 271833 125622 271838 125650
rect 271866 125622 295358 125650
rect 295386 125622 295391 125650
rect 271721 125566 271726 125594
rect 271754 125566 295470 125594
rect 295498 125566 295503 125594
rect 272113 124782 272118 124810
rect 272146 124782 276486 124810
rect 276514 124782 276519 124810
rect -480 124250 240 124348
rect -480 124236 28182 124250
rect 196 124222 28182 124236
rect 28210 124222 28215 124250
rect 297780 122514 298500 122612
rect 276985 122486 276990 122514
rect 277018 122500 298500 122514
rect 277018 122486 297836 122500
rect 196 117292 2366 117306
rect -480 117278 2366 117292
rect 2394 117278 2399 117306
rect -480 117180 240 117278
rect 295465 115990 295470 116018
rect 295498 116004 297836 116018
rect 295498 115990 298500 116004
rect 297780 115892 298500 115990
rect -480 110138 240 110236
rect -480 110124 28126 110138
rect 196 110110 28126 110124
rect 28154 110110 28159 110138
rect 297780 109284 298500 109396
rect 58697 107422 58702 107450
rect 58730 107422 75390 107450
rect 75418 107422 75423 107450
rect 57241 107366 57246 107394
rect 57274 107366 77742 107394
rect 77770 107366 77775 107394
rect 52985 107310 52990 107338
rect 53018 107310 74718 107338
rect 74746 107310 74751 107338
rect 47273 107254 47278 107282
rect 47306 107254 74046 107282
rect 74074 107254 74079 107282
rect 41561 107198 41566 107226
rect 41594 107198 73374 107226
rect 73402 107198 73407 107226
rect 35849 107142 35854 107170
rect 35882 107142 72702 107170
rect 72730 107142 72735 107170
rect 24425 107086 24430 107114
rect 24458 107086 71358 107114
rect 71386 107086 71391 107114
rect 43465 106638 43470 106666
rect 43498 106638 45150 106666
rect 45178 106638 45183 106666
rect 47161 106638 47166 106666
rect 47194 106638 49182 106666
rect 49210 106638 49215 106666
rect 64409 106638 64414 106666
rect 64442 106638 66766 106666
rect 66794 106638 66799 106666
rect 66873 106638 66878 106666
rect 66906 106638 68222 106666
rect 68250 106638 68255 106666
rect 78073 106638 78078 106666
rect 78106 106638 81550 106666
rect 81578 106638 81583 106666
rect 30137 106582 30142 106610
rect 30170 106582 37366 106610
rect 37394 106582 37399 106610
rect 39657 106582 39662 106610
rect 39690 106582 43806 106610
rect 43834 106582 43839 106610
rect 48281 106582 48286 106610
rect 48314 106582 51086 106610
rect 51114 106582 51119 106610
rect 51865 106582 51870 106610
rect 51898 106582 62510 106610
rect 62538 106582 62543 106610
rect 68441 106582 68446 106610
rect 68474 106582 73934 106610
rect 73962 106582 73967 106610
rect 32041 106526 32046 106554
rect 32074 106526 41118 106554
rect 41146 106526 41151 106554
rect 55225 106526 55230 106554
rect 55258 106526 72030 106554
rect 72058 106526 72063 106554
rect 78745 106526 78750 106554
rect 78778 106526 87262 106554
rect 87290 106526 87295 106554
rect 28233 106470 28238 106498
rect 28266 106470 39774 106498
rect 39802 106470 39807 106498
rect 57913 106470 57918 106498
rect 57946 106470 79646 106498
rect 79674 106470 79679 106498
rect 26329 106414 26334 106442
rect 26362 106414 39102 106442
rect 39130 106414 39135 106442
rect 53209 106414 53214 106442
rect 53242 106414 66318 106442
rect 66346 106414 66351 106442
rect 66985 106414 66990 106442
rect 67018 106414 91070 106442
rect 91098 106414 91103 106442
rect 22521 106358 22526 106386
rect 22554 106358 37758 106386
rect 37786 106358 37791 106386
rect 49961 106358 49966 106386
rect 49994 106358 54894 106386
rect 54922 106358 54927 106386
rect 59257 106358 59262 106386
rect 59290 106358 83454 106386
rect 83482 106358 83487 106386
rect 18713 106302 18718 106330
rect 18746 106302 34846 106330
rect 34874 106302 34879 106330
rect 49849 106302 49854 106330
rect 49882 106302 56798 106330
rect 56826 106302 56831 106330
rect 59929 106302 59934 106330
rect 59962 106302 85358 106330
rect 85386 106302 85391 106330
rect 20617 106246 20622 106274
rect 20650 106246 37086 106274
rect 37114 106246 37119 106274
rect 37753 106246 37758 106274
rect 37786 106246 43134 106274
rect 43162 106246 43167 106274
rect 51641 106246 51646 106274
rect 51674 106246 60606 106274
rect 60634 106246 60639 106274
rect 61273 106246 61278 106274
rect 61306 106246 89166 106274
rect 89194 106246 89199 106274
rect 196 103180 3150 103194
rect -480 103166 3150 103180
rect 3178 103166 3183 103194
rect -480 103068 240 103166
rect 297780 102690 298500 102788
rect 276929 102662 276934 102690
rect 276962 102676 298500 102690
rect 276962 102662 297836 102676
rect 295353 96166 295358 96194
rect 295386 96180 297836 96194
rect 295386 96166 298500 96180
rect -480 96026 240 96124
rect 297780 96068 298500 96166
rect -480 96012 6286 96026
rect 196 95998 6286 96012
rect 6314 95998 6319 96026
rect 297780 89460 298500 89572
rect -480 89026 240 89068
rect -480 88998 3990 89026
rect 4018 88998 4023 89026
rect -480 88956 240 88998
rect 297780 82866 298500 82964
rect 276873 82838 276878 82866
rect 276906 82852 298500 82866
rect 276906 82838 297836 82852
rect 196 82012 3934 82026
rect -480 81998 3934 82012
rect 3962 81998 3967 82026
rect -480 81900 240 81998
rect 295241 76342 295246 76370
rect 295274 76356 297836 76370
rect 295274 76342 298500 76356
rect 297780 76244 298500 76342
rect 19259 75334 19278 75362
rect 19306 75334 19311 75362
rect 19259 75110 19278 75138
rect 19306 75110 19311 75138
rect -480 74858 240 74956
rect -480 74844 7126 74858
rect 196 74830 7126 74844
rect 7154 74830 7159 74858
rect 18881 74718 18886 74746
rect 18914 74718 21406 74746
rect 21434 74718 21439 74746
rect 84457 73878 84462 73906
rect 84490 73878 90286 73906
rect 90314 73878 90319 73906
rect 82441 73822 82446 73850
rect 82474 73822 89502 73850
rect 89530 73822 89535 73850
rect 26441 73766 26446 73794
rect 26474 73766 32046 73794
rect 32074 73766 32079 73794
rect 88489 73766 88494 73794
rect 88522 73766 96166 73794
rect 96194 73766 96199 73794
rect 16137 73710 16142 73738
rect 16170 73710 25998 73738
rect 26026 73710 26031 73738
rect 29465 73710 29470 73738
rect 29498 73710 35406 73738
rect 35434 73710 35439 73738
rect 79081 73710 79086 73738
rect 79114 73710 88606 73738
rect 88634 73710 88639 73738
rect 14289 73654 14294 73682
rect 14322 73654 24654 73682
rect 24682 73654 24687 73682
rect 28569 73654 28574 73682
rect 28602 73654 34734 73682
rect 34762 73654 34767 73682
rect 87145 73654 87150 73682
rect 87178 73654 97846 73682
rect 97874 73654 97879 73682
rect 13281 73598 13286 73626
rect 13314 73598 23982 73626
rect 24010 73598 24015 73626
rect 24761 73598 24766 73626
rect 24794 73598 31374 73626
rect 31402 73598 31407 73626
rect 62281 73598 62286 73626
rect 62314 73598 65198 73626
rect 65226 73598 65231 73626
rect 66985 73598 66990 73626
rect 67018 73598 70966 73626
rect 70994 73598 70999 73626
rect 77065 73598 77070 73626
rect 77098 73598 87766 73626
rect 87794 73598 87799 73626
rect 89161 73598 89166 73626
rect 89194 73598 99526 73626
rect 99554 73598 99559 73626
rect 10425 73542 10430 73570
rect 10458 73542 21966 73570
rect 21994 73542 21999 73570
rect 23921 73542 23926 73570
rect 23954 73542 30702 73570
rect 30730 73542 30735 73570
rect 56905 73542 56910 73570
rect 56938 73542 59934 73570
rect 59962 73542 59967 73570
rect 74377 73542 74382 73570
rect 74410 73542 84686 73570
rect 84714 73542 84719 73570
rect 85129 73542 85134 73570
rect 85162 73542 96278 73570
rect 96306 73542 96311 73570
rect 9473 73486 9478 73514
rect 9506 73486 21294 73514
rect 21322 73486 21327 73514
rect 21849 73486 21854 73514
rect 21882 73486 30030 73514
rect 30058 73486 30063 73514
rect 30417 73486 30422 73514
rect 30450 73486 36078 73514
rect 36106 73486 36111 73514
rect 38985 73486 38990 73514
rect 39018 73486 42126 73514
rect 42154 73486 42159 73514
rect 62953 73486 62958 73514
rect 62986 73486 67774 73514
rect 67802 73486 67807 73514
rect 68329 73486 68334 73514
rect 68362 73486 72646 73514
rect 72674 73486 72679 73514
rect 81097 73486 81102 73514
rect 81130 73486 93646 73514
rect 93674 73486 93679 73514
rect 54217 73262 54222 73290
rect 54250 73262 56126 73290
rect 56154 73262 56159 73290
rect 54889 73206 54894 73234
rect 54922 73206 57134 73234
rect 57162 73206 57167 73234
rect 64969 73206 64974 73234
rect 65002 73206 69286 73234
rect 69314 73206 69319 73234
rect 24033 73150 24038 73178
rect 24066 73150 28686 73178
rect 28714 73150 28719 73178
rect 41841 73150 41846 73178
rect 41874 73150 44142 73178
rect 44170 73150 44175 73178
rect 52201 73150 52206 73178
rect 52234 73150 53270 73178
rect 53298 73150 53303 73178
rect 53545 73150 53550 73178
rect 53578 73150 55174 73178
rect 55202 73150 55207 73178
rect 66313 73150 66318 73178
rect 66346 73150 68446 73178
rect 68474 73150 68479 73178
rect 71017 73150 71022 73178
rect 71050 73150 73486 73178
rect 73514 73150 73519 73178
rect 18489 73094 18494 73122
rect 18522 73094 19278 73122
rect 19306 73094 19311 73122
rect 24873 73094 24878 73122
rect 24906 73094 29358 73122
rect 29386 73094 29391 73122
rect 34841 73094 34846 73122
rect 34874 73094 38766 73122
rect 38794 73094 38799 73122
rect 43745 73094 43750 73122
rect 43778 73094 45486 73122
rect 45514 73094 45519 73122
rect 51529 73094 51534 73122
rect 51562 73094 52318 73122
rect 52346 73094 52351 73122
rect 52873 73094 52878 73122
rect 52906 73094 54166 73122
rect 54194 73094 54199 73122
rect 58921 73094 58926 73122
rect 58954 73094 62790 73122
rect 62818 73094 62823 73122
rect 64297 73094 64302 73122
rect 64330 73094 65086 73122
rect 65114 73094 65119 73122
rect 65641 73094 65646 73122
rect 65674 73094 66766 73122
rect 66794 73094 66799 73122
rect 69001 73094 69006 73122
rect 69034 73094 72758 73122
rect 72786 73094 72791 73122
rect 73033 73094 73038 73122
rect 73066 73094 75166 73122
rect 75194 73094 75199 73122
rect 79753 73094 79758 73122
rect 79786 73094 80206 73122
rect 80234 73094 80239 73122
rect 297780 69636 298500 69748
rect 196 67900 2310 67914
rect -480 67886 2310 67900
rect 2338 67886 2343 67914
rect -480 67788 240 67886
rect 297780 63042 298500 63140
rect 276145 63014 276150 63042
rect 276178 63028 298500 63042
rect 276178 63014 297836 63028
rect 196 60844 3878 60858
rect -480 60830 3878 60844
rect 3906 60830 3911 60858
rect -480 60732 240 60830
rect 297780 56434 298500 56532
rect 276817 56406 276822 56434
rect 276850 56420 298500 56434
rect 276850 56406 297836 56420
rect -480 53746 240 53788
rect -480 53718 2254 53746
rect 2282 53718 2287 53746
rect -480 53676 240 53718
rect 297780 49812 298500 49924
rect 196 46732 2198 46746
rect -480 46718 2198 46732
rect 2226 46718 2231 46746
rect -480 46620 240 46718
rect 297780 43218 298500 43316
rect 276033 43190 276038 43218
rect 276066 43204 298500 43218
rect 276066 43190 297836 43204
rect 196 39676 3094 39690
rect -480 39662 3094 39676
rect 3122 39662 3127 39690
rect -480 39564 240 39662
rect 297780 36610 298500 36708
rect 276761 36582 276766 36610
rect 276794 36596 298500 36610
rect 276794 36582 297836 36596
rect 196 32620 3822 32634
rect -480 32606 3822 32620
rect 3850 32606 3855 32634
rect -480 32508 240 32606
rect 297780 29988 298500 30100
rect 196 25564 5446 25578
rect -480 25550 5446 25564
rect 5474 25550 5479 25578
rect -480 25452 240 25550
rect 297780 23394 298500 23492
rect 276089 23366 276094 23394
rect 276122 23380 298500 23394
rect 276122 23366 297836 23380
rect -480 18466 240 18508
rect -480 18438 3766 18466
rect 3794 18438 3799 18466
rect -480 18396 240 18438
rect 297780 16842 298500 16884
rect 275977 16814 275982 16842
rect 276010 16814 298500 16842
rect 297780 16772 298500 16814
rect 196 11452 2142 11466
rect -480 11438 2142 11452
rect 2170 11438 2175 11466
rect -480 11340 240 11438
rect 297780 10164 298500 10276
rect 7569 7126 7574 7154
rect 7602 7126 19950 7154
rect 19978 7126 19983 7154
rect 269369 7126 269374 7154
rect 269402 7126 278166 7154
rect 278194 7126 278199 7154
rect 260801 6398 260806 6426
rect 260834 6398 278222 6426
rect 278250 6398 278255 6426
rect 249377 6342 249382 6370
rect 249410 6342 277214 6370
rect 277242 6342 277247 6370
rect 243665 6286 243670 6314
rect 243698 6286 278278 6314
rect 278306 6286 278311 6314
rect 252345 4606 252350 4634
rect 252378 4606 278054 4634
rect 278082 4606 278087 4634
rect 196 4396 2086 4410
rect -480 4382 2086 4396
rect 2114 4382 2119 4410
rect -480 4284 240 4382
rect 255201 3822 255206 3850
rect 255234 3822 275646 3850
rect 275674 3822 275679 3850
rect 246633 3766 246638 3794
rect 246666 3766 278110 3794
rect 278138 3766 278143 3794
rect 297780 3570 298500 3668
rect 275921 3542 275926 3570
rect 275954 3556 298500 3570
rect 275954 3542 297836 3556
rect 75721 3318 75726 3346
rect 75754 3318 86590 3346
rect 86618 3318 86623 3346
rect 77737 3262 77742 3290
rect 77770 3262 89446 3290
rect 89474 3262 89479 3290
rect 69673 3206 69678 3234
rect 69706 3206 78022 3234
rect 78050 3206 78055 3234
rect 80201 3206 80206 3234
rect 80234 3206 92302 3234
rect 92330 3206 92335 3234
rect 18153 3150 18158 3178
rect 18186 3150 27342 3178
rect 27370 3150 27375 3178
rect 70345 3150 70350 3178
rect 70378 3150 78974 3178
rect 79002 3150 79007 3178
rect 80425 3150 80430 3178
rect 80458 3150 93254 3178
rect 93282 3150 93287 3178
rect 17201 3094 17206 3122
rect 17234 3094 26670 3122
rect 26698 3094 26703 3122
rect 71689 3094 71694 3122
rect 71722 3094 80878 3122
rect 80906 3094 80911 3122
rect 81769 3094 81774 3122
rect 81802 3094 95158 3122
rect 95186 3094 95191 3122
rect 15297 3038 15302 3066
rect 15330 3038 25326 3066
rect 25354 3038 25359 3066
rect 72361 3038 72366 3066
rect 72394 3038 81830 3066
rect 81858 3038 81863 3066
rect 83785 3038 83790 3066
rect 83818 3038 98014 3066
rect 98042 3038 98047 3066
rect 266625 3038 266630 3066
rect 266658 3038 276430 3066
rect 276458 3038 276463 3066
rect 12441 2982 12446 3010
rect 12474 2982 23310 3010
rect 23338 2982 23343 3010
rect 73705 2982 73710 3010
rect 73738 2982 83734 3010
rect 83762 2982 83767 3010
rect 85801 2982 85806 3010
rect 85834 2982 100870 3010
rect 100898 2982 100903 3010
rect 263713 2982 263718 3010
rect 263746 2982 276374 3010
rect 276402 2982 276407 3010
rect 8633 2926 8638 2954
rect 8666 2926 20622 2954
rect 20650 2926 20655 2954
rect 76393 2926 76398 2954
rect 76426 2926 87542 2954
rect 87570 2926 87575 2954
rect 87817 2926 87822 2954
rect 87850 2926 103726 2954
rect 103754 2926 103759 2954
rect 149305 2926 149310 2954
rect 149338 2926 157990 2954
rect 158018 2926 158023 2954
rect 258057 2926 258062 2954
rect 258090 2926 275590 2954
rect 275618 2926 275623 2954
rect 88601 2534 88606 2562
rect 88634 2534 91350 2562
rect 91378 2534 91383 2562
rect 37193 2478 37198 2506
rect 37226 2478 40782 2506
rect 40810 2478 40815 2506
rect 55561 2478 55566 2506
rect 55594 2478 58030 2506
rect 58058 2478 58063 2506
rect 59593 2478 59598 2506
rect 59626 2478 63742 2506
rect 63770 2478 63775 2506
rect 143817 2478 143822 2506
rect 143850 2478 145950 2506
rect 145978 2478 145983 2506
rect 277825 2478 277830 2506
rect 277858 2478 280798 2506
rect 280826 2478 280831 2506
rect 36241 2422 36246 2450
rect 36274 2422 40110 2450
rect 40138 2422 40143 2450
rect 44809 2422 44814 2450
rect 44842 2422 46158 2450
rect 46186 2422 46191 2450
rect 65081 2422 65086 2450
rect 65114 2422 70406 2450
rect 70434 2422 70439 2450
rect 72641 2422 72646 2450
rect 72674 2422 76118 2450
rect 76146 2422 76151 2450
rect 147961 2422 147966 2450
rect 147994 2422 152278 2450
rect 152306 2422 152311 2450
rect 20953 2366 20958 2394
rect 20986 2366 24878 2394
rect 24906 2366 24911 2394
rect 27706 2366 34062 2394
rect 34090 2366 34095 2394
rect 96273 2366 96278 2394
rect 96306 2366 99974 2394
rect 100002 2366 100007 2394
rect 22750 2254 24038 2282
rect 24066 2254 24071 2282
rect 27673 2254 27678 2282
rect 27706 2254 27734 2366
rect 32433 2310 32438 2338
rect 32466 2310 37422 2338
rect 37450 2310 37455 2338
rect 38145 2310 38150 2338
rect 38178 2310 41454 2338
rect 41482 2310 41487 2338
rect 68441 2310 68446 2338
rect 68474 2310 73262 2338
rect 73290 2310 73295 2338
rect 73481 2310 73486 2338
rect 73514 2310 79926 2338
rect 79954 2310 79959 2338
rect 89497 2310 89502 2338
rect 89530 2310 96110 2338
rect 96138 2310 96143 2338
rect 96217 2310 96222 2338
rect 96250 2310 97230 2338
rect 97258 2310 97263 2338
rect 97841 2310 97846 2338
rect 97874 2310 102774 2338
rect 102802 2310 102807 2338
rect 33385 2254 33390 2282
rect 33418 2254 38094 2282
rect 38122 2254 38127 2282
rect 60937 2254 60942 2282
rect 60970 2254 65646 2282
rect 65674 2254 65679 2282
rect 67657 2254 67662 2282
rect 67690 2254 75166 2282
rect 75194 2254 75199 2282
rect 90281 2254 90286 2282
rect 90314 2254 98966 2282
rect 98994 2254 98999 2282
rect 150649 2254 150654 2282
rect 150682 2254 163702 2282
rect 163730 2254 163735 2282
rect 11489 2198 11494 2226
rect 11522 2198 22638 2226
rect 22666 2198 22671 2226
rect 22750 2170 22778 2254
rect 24817 2198 24822 2226
rect 24850 2198 26446 2226
rect 26474 2198 26479 2226
rect 26721 2198 26726 2226
rect 26754 2198 33334 2226
rect 33362 2198 33367 2226
rect 56233 2198 56238 2226
rect 56266 2198 58982 2226
rect 59010 2198 59015 2226
rect 60265 2198 60270 2226
rect 60298 2198 64694 2226
rect 64722 2198 64727 2226
rect 72753 2198 72758 2226
rect 72786 2198 77070 2226
rect 77098 2198 77103 2226
rect 78409 2198 78414 2226
rect 78442 2198 90398 2226
rect 90426 2198 90431 2226
rect 92386 2198 97090 2226
rect 97225 2198 97230 2226
rect 97258 2198 104678 2226
rect 104706 2198 104711 2226
rect 151321 2198 151326 2226
rect 151354 2198 166558 2226
rect 166586 2198 166591 2226
rect 92386 2170 92414 2198
rect 97062 2170 97090 2198
rect 6673 2142 6678 2170
rect 6706 2142 18494 2170
rect 18522 2142 18527 2170
rect 20057 2142 20062 2170
rect 20090 2142 22778 2170
rect 22913 2142 22918 2170
rect 22946 2142 23926 2170
rect 23954 2142 23959 2170
rect 25769 2142 25774 2170
rect 25802 2142 32718 2170
rect 32746 2142 32751 2170
rect 34230 2142 36750 2170
rect 36778 2142 36783 2170
rect 41001 2142 41006 2170
rect 41034 2142 43470 2170
rect 43498 2142 43503 2170
rect 45761 2142 45766 2170
rect 45794 2142 46830 2170
rect 46858 2142 46863 2170
rect 61609 2142 61614 2170
rect 61642 2142 66598 2170
rect 66626 2142 66631 2170
rect 66761 2142 66766 2170
rect 66794 2142 72310 2170
rect 72338 2142 72343 2170
rect 75217 2142 75222 2170
rect 75250 2142 82782 2170
rect 82810 2142 82815 2170
rect 83113 2142 83118 2170
rect 83146 2142 92414 2170
rect 93641 2142 93646 2170
rect 93674 2142 94206 2170
rect 94234 2142 94239 2170
rect 97057 2142 97062 2170
rect 97090 2142 97095 2170
rect 99521 2142 99526 2170
rect 99554 2142 105630 2170
rect 105658 2142 105663 2170
rect 135193 2142 135198 2170
rect 135226 2142 143934 2170
rect 143962 2142 143967 2170
rect 151993 2142 151998 2170
rect 152026 2142 169414 2170
rect 169442 2142 169447 2170
rect 277713 2142 277718 2170
rect 277746 2142 283654 2170
rect 283682 2142 283687 2170
rect 34230 2114 34258 2142
rect 5777 2086 5782 2114
rect 5810 2086 18886 2114
rect 18914 2086 18919 2114
rect 19105 2086 19110 2114
rect 19138 2086 28014 2114
rect 28042 2086 28047 2114
rect 31481 2086 31486 2114
rect 31514 2086 34258 2114
rect 34337 2086 34342 2114
rect 34370 2086 34846 2114
rect 34874 2086 34879 2114
rect 35233 2086 35238 2114
rect 35266 2086 39438 2114
rect 39466 2086 39471 2114
rect 40049 2086 40054 2114
rect 40082 2086 42798 2114
rect 42826 2086 42831 2114
rect 42905 2086 42910 2114
rect 42938 2086 44758 2114
rect 44786 2086 44791 2114
rect 46713 2086 46718 2114
rect 46746 2086 47502 2114
rect 47530 2086 47535 2114
rect 47665 2086 47670 2114
rect 47698 2086 48174 2114
rect 48202 2086 48207 2114
rect 57577 2086 57582 2114
rect 57610 2086 60886 2114
rect 60914 2086 60919 2114
rect 65193 2086 65198 2114
rect 65226 2086 67550 2114
rect 67578 2086 67583 2114
rect 67769 2086 67774 2114
rect 67802 2086 68502 2114
rect 68530 2086 68535 2114
rect 68866 2086 69454 2114
rect 69482 2086 69487 2114
rect 70961 2086 70966 2114
rect 70994 2086 74214 2114
rect 74242 2086 74247 2114
rect 75049 2086 75054 2114
rect 75082 2086 85694 2114
rect 85722 2086 85727 2114
rect 86473 2086 86478 2114
rect 86506 2086 101822 2114
rect 101850 2086 101855 2114
rect 129537 2086 129542 2114
rect 129570 2086 142590 2114
rect 142618 2086 142623 2114
rect 147289 2086 147294 2114
rect 147322 2086 149422 2114
rect 149450 2086 149455 2114
rect 152665 2086 152670 2114
rect 152698 2086 172270 2114
rect 172298 2086 172303 2114
rect 272337 2086 272342 2114
rect 272370 2086 276486 2114
rect 276514 2086 276519 2114
rect 277601 2086 277606 2114
rect 277634 2086 286510 2114
rect 286538 2086 286543 2114
rect 68866 2058 68894 2086
rect 23865 2030 23870 2058
rect 23898 2030 24766 2058
rect 24794 2030 24799 2058
rect 58249 2030 58254 2058
rect 58282 2030 61838 2058
rect 61866 2030 61871 2058
rect 63625 2030 63630 2058
rect 63658 2030 68894 2058
rect 69281 2030 69286 2058
rect 69314 2030 71414 2058
rect 71442 2030 71447 2058
rect 87761 2030 87766 2058
rect 87794 2030 88494 2058
rect 88522 2030 88527 2058
rect 140961 2030 140966 2058
rect 140994 2030 145278 2058
rect 145306 2030 145311 2058
rect 159161 2030 159166 2058
rect 159194 2030 160846 2058
rect 160874 2030 160879 2058
<< via3 >>
rect 275926 294294 275954 294322
rect 3766 293566 3794 293594
rect 271726 287686 271754 287714
rect 2086 286510 2114 286538
rect 295246 281078 295274 281106
rect 5446 279454 5474 279482
rect 275086 274470 275114 274498
rect 3094 272398 3122 272426
rect 278446 267862 278474 267890
rect 2142 265342 2170 265370
rect 295302 261254 295330 261282
rect 5502 258286 5530 258314
rect 272566 254646 272594 254674
rect 3822 251230 3850 251258
rect 272622 248038 272650 248066
rect 2198 244174 2226 244202
rect 295358 241430 295386 241458
rect 5558 237118 5586 237146
rect 273406 234822 273434 234850
rect 3878 230062 3906 230090
rect 277606 228214 277634 228242
rect 2254 223006 2282 223034
rect 295414 221606 295442 221634
rect 5614 215950 5642 215978
rect 272678 215054 272706 215082
rect 3934 208894 3962 208922
rect 271782 208390 271810 208418
rect 6286 201838 6314 201866
rect 295470 201782 295498 201810
rect 276766 195174 276794 195202
rect 6342 194782 6370 194810
rect 271838 188566 271866 188594
rect 4942 187726 4970 187754
rect 272734 181958 272762 181986
rect 2310 180670 2338 180698
rect 271894 175350 271922 175378
rect 3150 173614 3178 173642
rect 271950 168742 271978 168770
rect 3990 166558 4018 166586
rect 272790 162134 272818 162162
rect 207046 162022 207074 162050
rect 207046 161742 207074 161770
rect 6398 159502 6426 159530
rect 275926 157654 275954 157682
rect 271726 157206 271754 157234
rect 295246 156758 295274 156786
rect 275086 156310 275114 156338
rect 3766 156086 3794 156114
rect 278446 155862 278474 155890
rect 2086 155526 2114 155554
rect 271726 155526 271754 155554
rect 295302 155414 295330 155442
rect 5446 154966 5474 154994
rect 272566 154966 272594 154994
rect 272622 154518 272650 154546
rect 3094 154406 3122 154434
rect 295358 154070 295386 154098
rect 2142 153846 2170 153874
rect 273406 153622 273434 153650
rect 5502 153286 5530 153314
rect 277606 153174 277634 153202
rect 3822 152726 3850 152754
rect 295414 152726 295442 152754
rect 2086 152446 2114 152474
rect 272678 152278 272706 152306
rect 2198 152166 2226 152194
rect 271782 151830 271810 151858
rect 5558 151606 5586 151634
rect 295470 151382 295498 151410
rect 3878 151046 3906 151074
rect 276766 150934 276794 150962
rect 2254 150486 2282 150514
rect 271838 150486 271866 150514
rect 272734 150038 272762 150066
rect 5614 149926 5642 149954
rect 271894 149590 271922 149618
rect 3934 149366 3962 149394
rect 271950 149142 271978 149170
rect 6286 148806 6314 148834
rect 272790 148694 272818 148722
rect 6342 148246 6370 148274
rect 271726 148246 271754 148274
rect 4942 147686 4970 147714
rect 271894 147350 271922 147378
rect 2310 147126 2338 147154
rect 271782 146902 271810 146930
rect 3150 146566 3178 146594
rect 3990 146006 4018 146034
rect 276990 146006 277018 146034
rect 271726 145558 271754 145586
rect 6398 145446 6426 145474
rect 2478 145390 2506 145418
rect 2086 144886 2114 144914
rect 276934 144662 276962 144690
rect 2478 144326 2506 144354
rect 271838 144214 271866 144242
rect 2086 143766 2114 143794
rect 276878 143318 276906 143346
rect 28238 143206 28266 143234
rect 271950 142870 271978 142898
rect 28182 142646 28210 142674
rect 271894 142310 271922 142338
rect 2366 142086 2394 142114
rect 276150 141974 276178 142002
rect 28126 141526 28154 141554
rect 276822 141526 276850 141554
rect 3150 140966 3178 140994
rect 276038 140630 276066 140658
rect 6286 140406 6314 140434
rect 276766 140182 276794 140210
rect 3990 139846 4018 139874
rect 3934 139286 3962 139314
rect 276094 139286 276122 139314
rect 275982 138838 276010 138866
rect 7126 138726 7154 138754
rect 2086 138446 2114 138474
rect 2310 138166 2338 138194
rect 275926 137942 275954 137970
rect 3878 137606 3906 137634
rect 2254 137046 2282 137074
rect 2198 136486 2226 136514
rect 3094 135926 3122 135954
rect 271782 135702 271810 135730
rect 3822 135366 3850 135394
rect 5446 134806 5474 134834
rect 3766 134246 3794 134274
rect 2142 133686 2170 133714
rect 2086 133126 2114 133154
rect 21406 132566 21434 132594
rect 19278 132006 19306 132034
rect 28238 131278 28266 131306
rect 107086 126686 107114 126714
rect 107086 126350 107114 126378
rect 271950 125678 271978 125706
rect 295246 125678 295274 125706
rect 271838 125622 271866 125650
rect 295358 125622 295386 125650
rect 271726 125566 271754 125594
rect 295470 125566 295498 125594
rect 28182 124222 28210 124250
rect 276990 122486 277018 122514
rect 2366 117278 2394 117306
rect 295470 115990 295498 116018
rect 28126 110110 28154 110138
rect 3150 103166 3178 103194
rect 276934 102662 276962 102690
rect 295358 96166 295386 96194
rect 6286 95998 6314 96026
rect 3990 88998 4018 89026
rect 276878 82838 276906 82866
rect 3934 81998 3962 82026
rect 295246 76342 295274 76370
rect 19278 75334 19306 75362
rect 19278 75110 19306 75138
rect 7126 74830 7154 74858
rect 21406 74718 21434 74746
rect 2310 67886 2338 67914
rect 276150 63014 276178 63042
rect 3878 60830 3906 60858
rect 276822 56406 276850 56434
rect 2254 53718 2282 53746
rect 2198 46718 2226 46746
rect 276038 43190 276066 43218
rect 3094 39662 3122 39690
rect 276766 36582 276794 36610
rect 3822 32606 3850 32634
rect 5446 25550 5474 25578
rect 276094 23366 276122 23394
rect 3766 18438 3794 18466
rect 275982 16814 276010 16842
rect 2142 11438 2170 11466
rect 2086 4382 2114 4410
rect 275926 3542 275954 3570
<< metal4 >>
rect -958 299086 -648 299134
rect -958 299058 -910 299086
rect -882 299058 -848 299086
rect -820 299058 -786 299086
rect -758 299058 -724 299086
rect -696 299058 -648 299086
rect -958 299024 -648 299058
rect -958 298996 -910 299024
rect -882 298996 -848 299024
rect -820 298996 -786 299024
rect -758 298996 -724 299024
rect -696 298996 -648 299024
rect -958 298962 -648 298996
rect -958 298934 -910 298962
rect -882 298934 -848 298962
rect -820 298934 -786 298962
rect -758 298934 -724 298962
rect -696 298934 -648 298962
rect -958 298900 -648 298934
rect -958 298872 -910 298900
rect -882 298872 -848 298900
rect -820 298872 -786 298900
rect -758 298872 -724 298900
rect -696 298872 -648 298900
rect -958 293175 -648 298872
rect -958 293147 -910 293175
rect -882 293147 -848 293175
rect -820 293147 -786 293175
rect -758 293147 -724 293175
rect -696 293147 -648 293175
rect -958 293113 -648 293147
rect -958 293085 -910 293113
rect -882 293085 -848 293113
rect -820 293085 -786 293113
rect -758 293085 -724 293113
rect -696 293085 -648 293113
rect -958 293051 -648 293085
rect -958 293023 -910 293051
rect -882 293023 -848 293051
rect -820 293023 -786 293051
rect -758 293023 -724 293051
rect -696 293023 -648 293051
rect -958 292989 -648 293023
rect -958 292961 -910 292989
rect -882 292961 -848 292989
rect -820 292961 -786 292989
rect -758 292961 -724 292989
rect -696 292961 -648 292989
rect -958 284175 -648 292961
rect -958 284147 -910 284175
rect -882 284147 -848 284175
rect -820 284147 -786 284175
rect -758 284147 -724 284175
rect -696 284147 -648 284175
rect -958 284113 -648 284147
rect -958 284085 -910 284113
rect -882 284085 -848 284113
rect -820 284085 -786 284113
rect -758 284085 -724 284113
rect -696 284085 -648 284113
rect -958 284051 -648 284085
rect -958 284023 -910 284051
rect -882 284023 -848 284051
rect -820 284023 -786 284051
rect -758 284023 -724 284051
rect -696 284023 -648 284051
rect -958 283989 -648 284023
rect -958 283961 -910 283989
rect -882 283961 -848 283989
rect -820 283961 -786 283989
rect -758 283961 -724 283989
rect -696 283961 -648 283989
rect -958 275175 -648 283961
rect -958 275147 -910 275175
rect -882 275147 -848 275175
rect -820 275147 -786 275175
rect -758 275147 -724 275175
rect -696 275147 -648 275175
rect -958 275113 -648 275147
rect -958 275085 -910 275113
rect -882 275085 -848 275113
rect -820 275085 -786 275113
rect -758 275085 -724 275113
rect -696 275085 -648 275113
rect -958 275051 -648 275085
rect -958 275023 -910 275051
rect -882 275023 -848 275051
rect -820 275023 -786 275051
rect -758 275023 -724 275051
rect -696 275023 -648 275051
rect -958 274989 -648 275023
rect -958 274961 -910 274989
rect -882 274961 -848 274989
rect -820 274961 -786 274989
rect -758 274961 -724 274989
rect -696 274961 -648 274989
rect -958 266175 -648 274961
rect -958 266147 -910 266175
rect -882 266147 -848 266175
rect -820 266147 -786 266175
rect -758 266147 -724 266175
rect -696 266147 -648 266175
rect -958 266113 -648 266147
rect -958 266085 -910 266113
rect -882 266085 -848 266113
rect -820 266085 -786 266113
rect -758 266085 -724 266113
rect -696 266085 -648 266113
rect -958 266051 -648 266085
rect -958 266023 -910 266051
rect -882 266023 -848 266051
rect -820 266023 -786 266051
rect -758 266023 -724 266051
rect -696 266023 -648 266051
rect -958 265989 -648 266023
rect -958 265961 -910 265989
rect -882 265961 -848 265989
rect -820 265961 -786 265989
rect -758 265961 -724 265989
rect -696 265961 -648 265989
rect -958 257175 -648 265961
rect -958 257147 -910 257175
rect -882 257147 -848 257175
rect -820 257147 -786 257175
rect -758 257147 -724 257175
rect -696 257147 -648 257175
rect -958 257113 -648 257147
rect -958 257085 -910 257113
rect -882 257085 -848 257113
rect -820 257085 -786 257113
rect -758 257085 -724 257113
rect -696 257085 -648 257113
rect -958 257051 -648 257085
rect -958 257023 -910 257051
rect -882 257023 -848 257051
rect -820 257023 -786 257051
rect -758 257023 -724 257051
rect -696 257023 -648 257051
rect -958 256989 -648 257023
rect -958 256961 -910 256989
rect -882 256961 -848 256989
rect -820 256961 -786 256989
rect -758 256961 -724 256989
rect -696 256961 -648 256989
rect -958 248175 -648 256961
rect -958 248147 -910 248175
rect -882 248147 -848 248175
rect -820 248147 -786 248175
rect -758 248147 -724 248175
rect -696 248147 -648 248175
rect -958 248113 -648 248147
rect -958 248085 -910 248113
rect -882 248085 -848 248113
rect -820 248085 -786 248113
rect -758 248085 -724 248113
rect -696 248085 -648 248113
rect -958 248051 -648 248085
rect -958 248023 -910 248051
rect -882 248023 -848 248051
rect -820 248023 -786 248051
rect -758 248023 -724 248051
rect -696 248023 -648 248051
rect -958 247989 -648 248023
rect -958 247961 -910 247989
rect -882 247961 -848 247989
rect -820 247961 -786 247989
rect -758 247961 -724 247989
rect -696 247961 -648 247989
rect -958 239175 -648 247961
rect -958 239147 -910 239175
rect -882 239147 -848 239175
rect -820 239147 -786 239175
rect -758 239147 -724 239175
rect -696 239147 -648 239175
rect -958 239113 -648 239147
rect -958 239085 -910 239113
rect -882 239085 -848 239113
rect -820 239085 -786 239113
rect -758 239085 -724 239113
rect -696 239085 -648 239113
rect -958 239051 -648 239085
rect -958 239023 -910 239051
rect -882 239023 -848 239051
rect -820 239023 -786 239051
rect -758 239023 -724 239051
rect -696 239023 -648 239051
rect -958 238989 -648 239023
rect -958 238961 -910 238989
rect -882 238961 -848 238989
rect -820 238961 -786 238989
rect -758 238961 -724 238989
rect -696 238961 -648 238989
rect -958 230175 -648 238961
rect -958 230147 -910 230175
rect -882 230147 -848 230175
rect -820 230147 -786 230175
rect -758 230147 -724 230175
rect -696 230147 -648 230175
rect -958 230113 -648 230147
rect -958 230085 -910 230113
rect -882 230085 -848 230113
rect -820 230085 -786 230113
rect -758 230085 -724 230113
rect -696 230085 -648 230113
rect -958 230051 -648 230085
rect -958 230023 -910 230051
rect -882 230023 -848 230051
rect -820 230023 -786 230051
rect -758 230023 -724 230051
rect -696 230023 -648 230051
rect -958 229989 -648 230023
rect -958 229961 -910 229989
rect -882 229961 -848 229989
rect -820 229961 -786 229989
rect -758 229961 -724 229989
rect -696 229961 -648 229989
rect -958 221175 -648 229961
rect -958 221147 -910 221175
rect -882 221147 -848 221175
rect -820 221147 -786 221175
rect -758 221147 -724 221175
rect -696 221147 -648 221175
rect -958 221113 -648 221147
rect -958 221085 -910 221113
rect -882 221085 -848 221113
rect -820 221085 -786 221113
rect -758 221085 -724 221113
rect -696 221085 -648 221113
rect -958 221051 -648 221085
rect -958 221023 -910 221051
rect -882 221023 -848 221051
rect -820 221023 -786 221051
rect -758 221023 -724 221051
rect -696 221023 -648 221051
rect -958 220989 -648 221023
rect -958 220961 -910 220989
rect -882 220961 -848 220989
rect -820 220961 -786 220989
rect -758 220961 -724 220989
rect -696 220961 -648 220989
rect -958 212175 -648 220961
rect -958 212147 -910 212175
rect -882 212147 -848 212175
rect -820 212147 -786 212175
rect -758 212147 -724 212175
rect -696 212147 -648 212175
rect -958 212113 -648 212147
rect -958 212085 -910 212113
rect -882 212085 -848 212113
rect -820 212085 -786 212113
rect -758 212085 -724 212113
rect -696 212085 -648 212113
rect -958 212051 -648 212085
rect -958 212023 -910 212051
rect -882 212023 -848 212051
rect -820 212023 -786 212051
rect -758 212023 -724 212051
rect -696 212023 -648 212051
rect -958 211989 -648 212023
rect -958 211961 -910 211989
rect -882 211961 -848 211989
rect -820 211961 -786 211989
rect -758 211961 -724 211989
rect -696 211961 -648 211989
rect -958 203175 -648 211961
rect -958 203147 -910 203175
rect -882 203147 -848 203175
rect -820 203147 -786 203175
rect -758 203147 -724 203175
rect -696 203147 -648 203175
rect -958 203113 -648 203147
rect -958 203085 -910 203113
rect -882 203085 -848 203113
rect -820 203085 -786 203113
rect -758 203085 -724 203113
rect -696 203085 -648 203113
rect -958 203051 -648 203085
rect -958 203023 -910 203051
rect -882 203023 -848 203051
rect -820 203023 -786 203051
rect -758 203023 -724 203051
rect -696 203023 -648 203051
rect -958 202989 -648 203023
rect -958 202961 -910 202989
rect -882 202961 -848 202989
rect -820 202961 -786 202989
rect -758 202961 -724 202989
rect -696 202961 -648 202989
rect -958 194175 -648 202961
rect -958 194147 -910 194175
rect -882 194147 -848 194175
rect -820 194147 -786 194175
rect -758 194147 -724 194175
rect -696 194147 -648 194175
rect -958 194113 -648 194147
rect -958 194085 -910 194113
rect -882 194085 -848 194113
rect -820 194085 -786 194113
rect -758 194085 -724 194113
rect -696 194085 -648 194113
rect -958 194051 -648 194085
rect -958 194023 -910 194051
rect -882 194023 -848 194051
rect -820 194023 -786 194051
rect -758 194023 -724 194051
rect -696 194023 -648 194051
rect -958 193989 -648 194023
rect -958 193961 -910 193989
rect -882 193961 -848 193989
rect -820 193961 -786 193989
rect -758 193961 -724 193989
rect -696 193961 -648 193989
rect -958 185175 -648 193961
rect -958 185147 -910 185175
rect -882 185147 -848 185175
rect -820 185147 -786 185175
rect -758 185147 -724 185175
rect -696 185147 -648 185175
rect -958 185113 -648 185147
rect -958 185085 -910 185113
rect -882 185085 -848 185113
rect -820 185085 -786 185113
rect -758 185085 -724 185113
rect -696 185085 -648 185113
rect -958 185051 -648 185085
rect -958 185023 -910 185051
rect -882 185023 -848 185051
rect -820 185023 -786 185051
rect -758 185023 -724 185051
rect -696 185023 -648 185051
rect -958 184989 -648 185023
rect -958 184961 -910 184989
rect -882 184961 -848 184989
rect -820 184961 -786 184989
rect -758 184961 -724 184989
rect -696 184961 -648 184989
rect -958 176175 -648 184961
rect -958 176147 -910 176175
rect -882 176147 -848 176175
rect -820 176147 -786 176175
rect -758 176147 -724 176175
rect -696 176147 -648 176175
rect -958 176113 -648 176147
rect -958 176085 -910 176113
rect -882 176085 -848 176113
rect -820 176085 -786 176113
rect -758 176085 -724 176113
rect -696 176085 -648 176113
rect -958 176051 -648 176085
rect -958 176023 -910 176051
rect -882 176023 -848 176051
rect -820 176023 -786 176051
rect -758 176023 -724 176051
rect -696 176023 -648 176051
rect -958 175989 -648 176023
rect -958 175961 -910 175989
rect -882 175961 -848 175989
rect -820 175961 -786 175989
rect -758 175961 -724 175989
rect -696 175961 -648 175989
rect -958 167175 -648 175961
rect -958 167147 -910 167175
rect -882 167147 -848 167175
rect -820 167147 -786 167175
rect -758 167147 -724 167175
rect -696 167147 -648 167175
rect -958 167113 -648 167147
rect -958 167085 -910 167113
rect -882 167085 -848 167113
rect -820 167085 -786 167113
rect -758 167085 -724 167113
rect -696 167085 -648 167113
rect -958 167051 -648 167085
rect -958 167023 -910 167051
rect -882 167023 -848 167051
rect -820 167023 -786 167051
rect -758 167023 -724 167051
rect -696 167023 -648 167051
rect -958 166989 -648 167023
rect -958 166961 -910 166989
rect -882 166961 -848 166989
rect -820 166961 -786 166989
rect -758 166961 -724 166989
rect -696 166961 -648 166989
rect -958 158175 -648 166961
rect -958 158147 -910 158175
rect -882 158147 -848 158175
rect -820 158147 -786 158175
rect -758 158147 -724 158175
rect -696 158147 -648 158175
rect -958 158113 -648 158147
rect -958 158085 -910 158113
rect -882 158085 -848 158113
rect -820 158085 -786 158113
rect -758 158085 -724 158113
rect -696 158085 -648 158113
rect -958 158051 -648 158085
rect -958 158023 -910 158051
rect -882 158023 -848 158051
rect -820 158023 -786 158051
rect -758 158023 -724 158051
rect -696 158023 -648 158051
rect -958 157989 -648 158023
rect -958 157961 -910 157989
rect -882 157961 -848 157989
rect -820 157961 -786 157989
rect -758 157961 -724 157989
rect -696 157961 -648 157989
rect -958 149175 -648 157961
rect -958 149147 -910 149175
rect -882 149147 -848 149175
rect -820 149147 -786 149175
rect -758 149147 -724 149175
rect -696 149147 -648 149175
rect -958 149113 -648 149147
rect -958 149085 -910 149113
rect -882 149085 -848 149113
rect -820 149085 -786 149113
rect -758 149085 -724 149113
rect -696 149085 -648 149113
rect -958 149051 -648 149085
rect -958 149023 -910 149051
rect -882 149023 -848 149051
rect -820 149023 -786 149051
rect -758 149023 -724 149051
rect -696 149023 -648 149051
rect -958 148989 -648 149023
rect -958 148961 -910 148989
rect -882 148961 -848 148989
rect -820 148961 -786 148989
rect -758 148961 -724 148989
rect -696 148961 -648 148989
rect -958 140175 -648 148961
rect -958 140147 -910 140175
rect -882 140147 -848 140175
rect -820 140147 -786 140175
rect -758 140147 -724 140175
rect -696 140147 -648 140175
rect -958 140113 -648 140147
rect -958 140085 -910 140113
rect -882 140085 -848 140113
rect -820 140085 -786 140113
rect -758 140085 -724 140113
rect -696 140085 -648 140113
rect -958 140051 -648 140085
rect -958 140023 -910 140051
rect -882 140023 -848 140051
rect -820 140023 -786 140051
rect -758 140023 -724 140051
rect -696 140023 -648 140051
rect -958 139989 -648 140023
rect -958 139961 -910 139989
rect -882 139961 -848 139989
rect -820 139961 -786 139989
rect -758 139961 -724 139989
rect -696 139961 -648 139989
rect -958 131175 -648 139961
rect -958 131147 -910 131175
rect -882 131147 -848 131175
rect -820 131147 -786 131175
rect -758 131147 -724 131175
rect -696 131147 -648 131175
rect -958 131113 -648 131147
rect -958 131085 -910 131113
rect -882 131085 -848 131113
rect -820 131085 -786 131113
rect -758 131085 -724 131113
rect -696 131085 -648 131113
rect -958 131051 -648 131085
rect -958 131023 -910 131051
rect -882 131023 -848 131051
rect -820 131023 -786 131051
rect -758 131023 -724 131051
rect -696 131023 -648 131051
rect -958 130989 -648 131023
rect -958 130961 -910 130989
rect -882 130961 -848 130989
rect -820 130961 -786 130989
rect -758 130961 -724 130989
rect -696 130961 -648 130989
rect -958 122175 -648 130961
rect -958 122147 -910 122175
rect -882 122147 -848 122175
rect -820 122147 -786 122175
rect -758 122147 -724 122175
rect -696 122147 -648 122175
rect -958 122113 -648 122147
rect -958 122085 -910 122113
rect -882 122085 -848 122113
rect -820 122085 -786 122113
rect -758 122085 -724 122113
rect -696 122085 -648 122113
rect -958 122051 -648 122085
rect -958 122023 -910 122051
rect -882 122023 -848 122051
rect -820 122023 -786 122051
rect -758 122023 -724 122051
rect -696 122023 -648 122051
rect -958 121989 -648 122023
rect -958 121961 -910 121989
rect -882 121961 -848 121989
rect -820 121961 -786 121989
rect -758 121961 -724 121989
rect -696 121961 -648 121989
rect -958 113175 -648 121961
rect -958 113147 -910 113175
rect -882 113147 -848 113175
rect -820 113147 -786 113175
rect -758 113147 -724 113175
rect -696 113147 -648 113175
rect -958 113113 -648 113147
rect -958 113085 -910 113113
rect -882 113085 -848 113113
rect -820 113085 -786 113113
rect -758 113085 -724 113113
rect -696 113085 -648 113113
rect -958 113051 -648 113085
rect -958 113023 -910 113051
rect -882 113023 -848 113051
rect -820 113023 -786 113051
rect -758 113023 -724 113051
rect -696 113023 -648 113051
rect -958 112989 -648 113023
rect -958 112961 -910 112989
rect -882 112961 -848 112989
rect -820 112961 -786 112989
rect -758 112961 -724 112989
rect -696 112961 -648 112989
rect -958 104175 -648 112961
rect -958 104147 -910 104175
rect -882 104147 -848 104175
rect -820 104147 -786 104175
rect -758 104147 -724 104175
rect -696 104147 -648 104175
rect -958 104113 -648 104147
rect -958 104085 -910 104113
rect -882 104085 -848 104113
rect -820 104085 -786 104113
rect -758 104085 -724 104113
rect -696 104085 -648 104113
rect -958 104051 -648 104085
rect -958 104023 -910 104051
rect -882 104023 -848 104051
rect -820 104023 -786 104051
rect -758 104023 -724 104051
rect -696 104023 -648 104051
rect -958 103989 -648 104023
rect -958 103961 -910 103989
rect -882 103961 -848 103989
rect -820 103961 -786 103989
rect -758 103961 -724 103989
rect -696 103961 -648 103989
rect -958 95175 -648 103961
rect -958 95147 -910 95175
rect -882 95147 -848 95175
rect -820 95147 -786 95175
rect -758 95147 -724 95175
rect -696 95147 -648 95175
rect -958 95113 -648 95147
rect -958 95085 -910 95113
rect -882 95085 -848 95113
rect -820 95085 -786 95113
rect -758 95085 -724 95113
rect -696 95085 -648 95113
rect -958 95051 -648 95085
rect -958 95023 -910 95051
rect -882 95023 -848 95051
rect -820 95023 -786 95051
rect -758 95023 -724 95051
rect -696 95023 -648 95051
rect -958 94989 -648 95023
rect -958 94961 -910 94989
rect -882 94961 -848 94989
rect -820 94961 -786 94989
rect -758 94961 -724 94989
rect -696 94961 -648 94989
rect -958 86175 -648 94961
rect -958 86147 -910 86175
rect -882 86147 -848 86175
rect -820 86147 -786 86175
rect -758 86147 -724 86175
rect -696 86147 -648 86175
rect -958 86113 -648 86147
rect -958 86085 -910 86113
rect -882 86085 -848 86113
rect -820 86085 -786 86113
rect -758 86085 -724 86113
rect -696 86085 -648 86113
rect -958 86051 -648 86085
rect -958 86023 -910 86051
rect -882 86023 -848 86051
rect -820 86023 -786 86051
rect -758 86023 -724 86051
rect -696 86023 -648 86051
rect -958 85989 -648 86023
rect -958 85961 -910 85989
rect -882 85961 -848 85989
rect -820 85961 -786 85989
rect -758 85961 -724 85989
rect -696 85961 -648 85989
rect -958 77175 -648 85961
rect -958 77147 -910 77175
rect -882 77147 -848 77175
rect -820 77147 -786 77175
rect -758 77147 -724 77175
rect -696 77147 -648 77175
rect -958 77113 -648 77147
rect -958 77085 -910 77113
rect -882 77085 -848 77113
rect -820 77085 -786 77113
rect -758 77085 -724 77113
rect -696 77085 -648 77113
rect -958 77051 -648 77085
rect -958 77023 -910 77051
rect -882 77023 -848 77051
rect -820 77023 -786 77051
rect -758 77023 -724 77051
rect -696 77023 -648 77051
rect -958 76989 -648 77023
rect -958 76961 -910 76989
rect -882 76961 -848 76989
rect -820 76961 -786 76989
rect -758 76961 -724 76989
rect -696 76961 -648 76989
rect -958 68175 -648 76961
rect -958 68147 -910 68175
rect -882 68147 -848 68175
rect -820 68147 -786 68175
rect -758 68147 -724 68175
rect -696 68147 -648 68175
rect -958 68113 -648 68147
rect -958 68085 -910 68113
rect -882 68085 -848 68113
rect -820 68085 -786 68113
rect -758 68085 -724 68113
rect -696 68085 -648 68113
rect -958 68051 -648 68085
rect -958 68023 -910 68051
rect -882 68023 -848 68051
rect -820 68023 -786 68051
rect -758 68023 -724 68051
rect -696 68023 -648 68051
rect -958 67989 -648 68023
rect -958 67961 -910 67989
rect -882 67961 -848 67989
rect -820 67961 -786 67989
rect -758 67961 -724 67989
rect -696 67961 -648 67989
rect -958 59175 -648 67961
rect -958 59147 -910 59175
rect -882 59147 -848 59175
rect -820 59147 -786 59175
rect -758 59147 -724 59175
rect -696 59147 -648 59175
rect -958 59113 -648 59147
rect -958 59085 -910 59113
rect -882 59085 -848 59113
rect -820 59085 -786 59113
rect -758 59085 -724 59113
rect -696 59085 -648 59113
rect -958 59051 -648 59085
rect -958 59023 -910 59051
rect -882 59023 -848 59051
rect -820 59023 -786 59051
rect -758 59023 -724 59051
rect -696 59023 -648 59051
rect -958 58989 -648 59023
rect -958 58961 -910 58989
rect -882 58961 -848 58989
rect -820 58961 -786 58989
rect -758 58961 -724 58989
rect -696 58961 -648 58989
rect -958 50175 -648 58961
rect -958 50147 -910 50175
rect -882 50147 -848 50175
rect -820 50147 -786 50175
rect -758 50147 -724 50175
rect -696 50147 -648 50175
rect -958 50113 -648 50147
rect -958 50085 -910 50113
rect -882 50085 -848 50113
rect -820 50085 -786 50113
rect -758 50085 -724 50113
rect -696 50085 -648 50113
rect -958 50051 -648 50085
rect -958 50023 -910 50051
rect -882 50023 -848 50051
rect -820 50023 -786 50051
rect -758 50023 -724 50051
rect -696 50023 -648 50051
rect -958 49989 -648 50023
rect -958 49961 -910 49989
rect -882 49961 -848 49989
rect -820 49961 -786 49989
rect -758 49961 -724 49989
rect -696 49961 -648 49989
rect -958 41175 -648 49961
rect -958 41147 -910 41175
rect -882 41147 -848 41175
rect -820 41147 -786 41175
rect -758 41147 -724 41175
rect -696 41147 -648 41175
rect -958 41113 -648 41147
rect -958 41085 -910 41113
rect -882 41085 -848 41113
rect -820 41085 -786 41113
rect -758 41085 -724 41113
rect -696 41085 -648 41113
rect -958 41051 -648 41085
rect -958 41023 -910 41051
rect -882 41023 -848 41051
rect -820 41023 -786 41051
rect -758 41023 -724 41051
rect -696 41023 -648 41051
rect -958 40989 -648 41023
rect -958 40961 -910 40989
rect -882 40961 -848 40989
rect -820 40961 -786 40989
rect -758 40961 -724 40989
rect -696 40961 -648 40989
rect -958 32175 -648 40961
rect -958 32147 -910 32175
rect -882 32147 -848 32175
rect -820 32147 -786 32175
rect -758 32147 -724 32175
rect -696 32147 -648 32175
rect -958 32113 -648 32147
rect -958 32085 -910 32113
rect -882 32085 -848 32113
rect -820 32085 -786 32113
rect -758 32085 -724 32113
rect -696 32085 -648 32113
rect -958 32051 -648 32085
rect -958 32023 -910 32051
rect -882 32023 -848 32051
rect -820 32023 -786 32051
rect -758 32023 -724 32051
rect -696 32023 -648 32051
rect -958 31989 -648 32023
rect -958 31961 -910 31989
rect -882 31961 -848 31989
rect -820 31961 -786 31989
rect -758 31961 -724 31989
rect -696 31961 -648 31989
rect -958 23175 -648 31961
rect -958 23147 -910 23175
rect -882 23147 -848 23175
rect -820 23147 -786 23175
rect -758 23147 -724 23175
rect -696 23147 -648 23175
rect -958 23113 -648 23147
rect -958 23085 -910 23113
rect -882 23085 -848 23113
rect -820 23085 -786 23113
rect -758 23085 -724 23113
rect -696 23085 -648 23113
rect -958 23051 -648 23085
rect -958 23023 -910 23051
rect -882 23023 -848 23051
rect -820 23023 -786 23051
rect -758 23023 -724 23051
rect -696 23023 -648 23051
rect -958 22989 -648 23023
rect -958 22961 -910 22989
rect -882 22961 -848 22989
rect -820 22961 -786 22989
rect -758 22961 -724 22989
rect -696 22961 -648 22989
rect -958 14175 -648 22961
rect -958 14147 -910 14175
rect -882 14147 -848 14175
rect -820 14147 -786 14175
rect -758 14147 -724 14175
rect -696 14147 -648 14175
rect -958 14113 -648 14147
rect -958 14085 -910 14113
rect -882 14085 -848 14113
rect -820 14085 -786 14113
rect -758 14085 -724 14113
rect -696 14085 -648 14113
rect -958 14051 -648 14085
rect -958 14023 -910 14051
rect -882 14023 -848 14051
rect -820 14023 -786 14051
rect -758 14023 -724 14051
rect -696 14023 -648 14051
rect -958 13989 -648 14023
rect -958 13961 -910 13989
rect -882 13961 -848 13989
rect -820 13961 -786 13989
rect -758 13961 -724 13989
rect -696 13961 -648 13989
rect -958 5175 -648 13961
rect -958 5147 -910 5175
rect -882 5147 -848 5175
rect -820 5147 -786 5175
rect -758 5147 -724 5175
rect -696 5147 -648 5175
rect -958 5113 -648 5147
rect -958 5085 -910 5113
rect -882 5085 -848 5113
rect -820 5085 -786 5113
rect -758 5085 -724 5113
rect -696 5085 -648 5113
rect -958 5051 -648 5085
rect -958 5023 -910 5051
rect -882 5023 -848 5051
rect -820 5023 -786 5051
rect -758 5023 -724 5051
rect -696 5023 -648 5051
rect -958 4989 -648 5023
rect -958 4961 -910 4989
rect -882 4961 -848 4989
rect -820 4961 -786 4989
rect -758 4961 -724 4989
rect -696 4961 -648 4989
rect -958 -560 -648 4961
rect -478 298606 -168 298654
rect -478 298578 -430 298606
rect -402 298578 -368 298606
rect -340 298578 -306 298606
rect -278 298578 -244 298606
rect -216 298578 -168 298606
rect -478 298544 -168 298578
rect -478 298516 -430 298544
rect -402 298516 -368 298544
rect -340 298516 -306 298544
rect -278 298516 -244 298544
rect -216 298516 -168 298544
rect -478 298482 -168 298516
rect -478 298454 -430 298482
rect -402 298454 -368 298482
rect -340 298454 -306 298482
rect -278 298454 -244 298482
rect -216 298454 -168 298482
rect -478 298420 -168 298454
rect -478 298392 -430 298420
rect -402 298392 -368 298420
rect -340 298392 -306 298420
rect -278 298392 -244 298420
rect -216 298392 -168 298420
rect -478 290175 -168 298392
rect -478 290147 -430 290175
rect -402 290147 -368 290175
rect -340 290147 -306 290175
rect -278 290147 -244 290175
rect -216 290147 -168 290175
rect -478 290113 -168 290147
rect -478 290085 -430 290113
rect -402 290085 -368 290113
rect -340 290085 -306 290113
rect -278 290085 -244 290113
rect -216 290085 -168 290113
rect -478 290051 -168 290085
rect -478 290023 -430 290051
rect -402 290023 -368 290051
rect -340 290023 -306 290051
rect -278 290023 -244 290051
rect -216 290023 -168 290051
rect -478 289989 -168 290023
rect -478 289961 -430 289989
rect -402 289961 -368 289989
rect -340 289961 -306 289989
rect -278 289961 -244 289989
rect -216 289961 -168 289989
rect -478 281175 -168 289961
rect 2709 298606 3019 299134
rect 2709 298578 2757 298606
rect 2785 298578 2819 298606
rect 2847 298578 2881 298606
rect 2909 298578 2943 298606
rect 2971 298578 3019 298606
rect 2709 298544 3019 298578
rect 2709 298516 2757 298544
rect 2785 298516 2819 298544
rect 2847 298516 2881 298544
rect 2909 298516 2943 298544
rect 2971 298516 3019 298544
rect 2709 298482 3019 298516
rect 2709 298454 2757 298482
rect 2785 298454 2819 298482
rect 2847 298454 2881 298482
rect 2909 298454 2943 298482
rect 2971 298454 3019 298482
rect 2709 298420 3019 298454
rect 2709 298392 2757 298420
rect 2785 298392 2819 298420
rect 2847 298392 2881 298420
rect 2909 298392 2943 298420
rect 2971 298392 3019 298420
rect 2709 290175 3019 298392
rect 4569 299086 4879 299134
rect 4569 299058 4617 299086
rect 4645 299058 4679 299086
rect 4707 299058 4741 299086
rect 4769 299058 4803 299086
rect 4831 299058 4879 299086
rect 4569 299024 4879 299058
rect 4569 298996 4617 299024
rect 4645 298996 4679 299024
rect 4707 298996 4741 299024
rect 4769 298996 4803 299024
rect 4831 298996 4879 299024
rect 4569 298962 4879 298996
rect 4569 298934 4617 298962
rect 4645 298934 4679 298962
rect 4707 298934 4741 298962
rect 4769 298934 4803 298962
rect 4831 298934 4879 298962
rect 4569 298900 4879 298934
rect 4569 298872 4617 298900
rect 4645 298872 4679 298900
rect 4707 298872 4741 298900
rect 4769 298872 4803 298900
rect 4831 298872 4879 298900
rect 2709 290147 2757 290175
rect 2785 290147 2819 290175
rect 2847 290147 2881 290175
rect 2909 290147 2943 290175
rect 2971 290147 3019 290175
rect 2709 290113 3019 290147
rect 2709 290085 2757 290113
rect 2785 290085 2819 290113
rect 2847 290085 2881 290113
rect 2909 290085 2943 290113
rect 2971 290085 3019 290113
rect 2709 290051 3019 290085
rect 2709 290023 2757 290051
rect 2785 290023 2819 290051
rect 2847 290023 2881 290051
rect 2909 290023 2943 290051
rect 2971 290023 3019 290051
rect 2709 289989 3019 290023
rect 2709 289961 2757 289989
rect 2785 289961 2819 289989
rect 2847 289961 2881 289989
rect 2909 289961 2943 289989
rect 2971 289961 3019 289989
rect -478 281147 -430 281175
rect -402 281147 -368 281175
rect -340 281147 -306 281175
rect -278 281147 -244 281175
rect -216 281147 -168 281175
rect -478 281113 -168 281147
rect -478 281085 -430 281113
rect -402 281085 -368 281113
rect -340 281085 -306 281113
rect -278 281085 -244 281113
rect -216 281085 -168 281113
rect -478 281051 -168 281085
rect -478 281023 -430 281051
rect -402 281023 -368 281051
rect -340 281023 -306 281051
rect -278 281023 -244 281051
rect -216 281023 -168 281051
rect -478 280989 -168 281023
rect -478 280961 -430 280989
rect -402 280961 -368 280989
rect -340 280961 -306 280989
rect -278 280961 -244 280989
rect -216 280961 -168 280989
rect -478 272175 -168 280961
rect -478 272147 -430 272175
rect -402 272147 -368 272175
rect -340 272147 -306 272175
rect -278 272147 -244 272175
rect -216 272147 -168 272175
rect -478 272113 -168 272147
rect -478 272085 -430 272113
rect -402 272085 -368 272113
rect -340 272085 -306 272113
rect -278 272085 -244 272113
rect -216 272085 -168 272113
rect -478 272051 -168 272085
rect -478 272023 -430 272051
rect -402 272023 -368 272051
rect -340 272023 -306 272051
rect -278 272023 -244 272051
rect -216 272023 -168 272051
rect -478 271989 -168 272023
rect -478 271961 -430 271989
rect -402 271961 -368 271989
rect -340 271961 -306 271989
rect -278 271961 -244 271989
rect -216 271961 -168 271989
rect -478 263175 -168 271961
rect -478 263147 -430 263175
rect -402 263147 -368 263175
rect -340 263147 -306 263175
rect -278 263147 -244 263175
rect -216 263147 -168 263175
rect -478 263113 -168 263147
rect -478 263085 -430 263113
rect -402 263085 -368 263113
rect -340 263085 -306 263113
rect -278 263085 -244 263113
rect -216 263085 -168 263113
rect -478 263051 -168 263085
rect -478 263023 -430 263051
rect -402 263023 -368 263051
rect -340 263023 -306 263051
rect -278 263023 -244 263051
rect -216 263023 -168 263051
rect -478 262989 -168 263023
rect -478 262961 -430 262989
rect -402 262961 -368 262989
rect -340 262961 -306 262989
rect -278 262961 -244 262989
rect -216 262961 -168 262989
rect -478 254175 -168 262961
rect -478 254147 -430 254175
rect -402 254147 -368 254175
rect -340 254147 -306 254175
rect -278 254147 -244 254175
rect -216 254147 -168 254175
rect -478 254113 -168 254147
rect -478 254085 -430 254113
rect -402 254085 -368 254113
rect -340 254085 -306 254113
rect -278 254085 -244 254113
rect -216 254085 -168 254113
rect -478 254051 -168 254085
rect -478 254023 -430 254051
rect -402 254023 -368 254051
rect -340 254023 -306 254051
rect -278 254023 -244 254051
rect -216 254023 -168 254051
rect -478 253989 -168 254023
rect -478 253961 -430 253989
rect -402 253961 -368 253989
rect -340 253961 -306 253989
rect -278 253961 -244 253989
rect -216 253961 -168 253989
rect -478 245175 -168 253961
rect -478 245147 -430 245175
rect -402 245147 -368 245175
rect -340 245147 -306 245175
rect -278 245147 -244 245175
rect -216 245147 -168 245175
rect -478 245113 -168 245147
rect -478 245085 -430 245113
rect -402 245085 -368 245113
rect -340 245085 -306 245113
rect -278 245085 -244 245113
rect -216 245085 -168 245113
rect -478 245051 -168 245085
rect -478 245023 -430 245051
rect -402 245023 -368 245051
rect -340 245023 -306 245051
rect -278 245023 -244 245051
rect -216 245023 -168 245051
rect -478 244989 -168 245023
rect -478 244961 -430 244989
rect -402 244961 -368 244989
rect -340 244961 -306 244989
rect -278 244961 -244 244989
rect -216 244961 -168 244989
rect -478 236175 -168 244961
rect -478 236147 -430 236175
rect -402 236147 -368 236175
rect -340 236147 -306 236175
rect -278 236147 -244 236175
rect -216 236147 -168 236175
rect -478 236113 -168 236147
rect -478 236085 -430 236113
rect -402 236085 -368 236113
rect -340 236085 -306 236113
rect -278 236085 -244 236113
rect -216 236085 -168 236113
rect -478 236051 -168 236085
rect -478 236023 -430 236051
rect -402 236023 -368 236051
rect -340 236023 -306 236051
rect -278 236023 -244 236051
rect -216 236023 -168 236051
rect -478 235989 -168 236023
rect -478 235961 -430 235989
rect -402 235961 -368 235989
rect -340 235961 -306 235989
rect -278 235961 -244 235989
rect -216 235961 -168 235989
rect -478 227175 -168 235961
rect -478 227147 -430 227175
rect -402 227147 -368 227175
rect -340 227147 -306 227175
rect -278 227147 -244 227175
rect -216 227147 -168 227175
rect -478 227113 -168 227147
rect -478 227085 -430 227113
rect -402 227085 -368 227113
rect -340 227085 -306 227113
rect -278 227085 -244 227113
rect -216 227085 -168 227113
rect -478 227051 -168 227085
rect -478 227023 -430 227051
rect -402 227023 -368 227051
rect -340 227023 -306 227051
rect -278 227023 -244 227051
rect -216 227023 -168 227051
rect -478 226989 -168 227023
rect -478 226961 -430 226989
rect -402 226961 -368 226989
rect -340 226961 -306 226989
rect -278 226961 -244 226989
rect -216 226961 -168 226989
rect -478 218175 -168 226961
rect -478 218147 -430 218175
rect -402 218147 -368 218175
rect -340 218147 -306 218175
rect -278 218147 -244 218175
rect -216 218147 -168 218175
rect -478 218113 -168 218147
rect -478 218085 -430 218113
rect -402 218085 -368 218113
rect -340 218085 -306 218113
rect -278 218085 -244 218113
rect -216 218085 -168 218113
rect -478 218051 -168 218085
rect -478 218023 -430 218051
rect -402 218023 -368 218051
rect -340 218023 -306 218051
rect -278 218023 -244 218051
rect -216 218023 -168 218051
rect -478 217989 -168 218023
rect -478 217961 -430 217989
rect -402 217961 -368 217989
rect -340 217961 -306 217989
rect -278 217961 -244 217989
rect -216 217961 -168 217989
rect -478 209175 -168 217961
rect -478 209147 -430 209175
rect -402 209147 -368 209175
rect -340 209147 -306 209175
rect -278 209147 -244 209175
rect -216 209147 -168 209175
rect -478 209113 -168 209147
rect -478 209085 -430 209113
rect -402 209085 -368 209113
rect -340 209085 -306 209113
rect -278 209085 -244 209113
rect -216 209085 -168 209113
rect -478 209051 -168 209085
rect -478 209023 -430 209051
rect -402 209023 -368 209051
rect -340 209023 -306 209051
rect -278 209023 -244 209051
rect -216 209023 -168 209051
rect -478 208989 -168 209023
rect -478 208961 -430 208989
rect -402 208961 -368 208989
rect -340 208961 -306 208989
rect -278 208961 -244 208989
rect -216 208961 -168 208989
rect -478 200175 -168 208961
rect -478 200147 -430 200175
rect -402 200147 -368 200175
rect -340 200147 -306 200175
rect -278 200147 -244 200175
rect -216 200147 -168 200175
rect -478 200113 -168 200147
rect -478 200085 -430 200113
rect -402 200085 -368 200113
rect -340 200085 -306 200113
rect -278 200085 -244 200113
rect -216 200085 -168 200113
rect -478 200051 -168 200085
rect -478 200023 -430 200051
rect -402 200023 -368 200051
rect -340 200023 -306 200051
rect -278 200023 -244 200051
rect -216 200023 -168 200051
rect -478 199989 -168 200023
rect -478 199961 -430 199989
rect -402 199961 -368 199989
rect -340 199961 -306 199989
rect -278 199961 -244 199989
rect -216 199961 -168 199989
rect -478 191175 -168 199961
rect -478 191147 -430 191175
rect -402 191147 -368 191175
rect -340 191147 -306 191175
rect -278 191147 -244 191175
rect -216 191147 -168 191175
rect -478 191113 -168 191147
rect -478 191085 -430 191113
rect -402 191085 -368 191113
rect -340 191085 -306 191113
rect -278 191085 -244 191113
rect -216 191085 -168 191113
rect -478 191051 -168 191085
rect -478 191023 -430 191051
rect -402 191023 -368 191051
rect -340 191023 -306 191051
rect -278 191023 -244 191051
rect -216 191023 -168 191051
rect -478 190989 -168 191023
rect -478 190961 -430 190989
rect -402 190961 -368 190989
rect -340 190961 -306 190989
rect -278 190961 -244 190989
rect -216 190961 -168 190989
rect -478 182175 -168 190961
rect -478 182147 -430 182175
rect -402 182147 -368 182175
rect -340 182147 -306 182175
rect -278 182147 -244 182175
rect -216 182147 -168 182175
rect -478 182113 -168 182147
rect -478 182085 -430 182113
rect -402 182085 -368 182113
rect -340 182085 -306 182113
rect -278 182085 -244 182113
rect -216 182085 -168 182113
rect -478 182051 -168 182085
rect -478 182023 -430 182051
rect -402 182023 -368 182051
rect -340 182023 -306 182051
rect -278 182023 -244 182051
rect -216 182023 -168 182051
rect -478 181989 -168 182023
rect -478 181961 -430 181989
rect -402 181961 -368 181989
rect -340 181961 -306 181989
rect -278 181961 -244 181989
rect -216 181961 -168 181989
rect -478 173175 -168 181961
rect -478 173147 -430 173175
rect -402 173147 -368 173175
rect -340 173147 -306 173175
rect -278 173147 -244 173175
rect -216 173147 -168 173175
rect -478 173113 -168 173147
rect -478 173085 -430 173113
rect -402 173085 -368 173113
rect -340 173085 -306 173113
rect -278 173085 -244 173113
rect -216 173085 -168 173113
rect -478 173051 -168 173085
rect -478 173023 -430 173051
rect -402 173023 -368 173051
rect -340 173023 -306 173051
rect -278 173023 -244 173051
rect -216 173023 -168 173051
rect -478 172989 -168 173023
rect -478 172961 -430 172989
rect -402 172961 -368 172989
rect -340 172961 -306 172989
rect -278 172961 -244 172989
rect -216 172961 -168 172989
rect -478 164175 -168 172961
rect -478 164147 -430 164175
rect -402 164147 -368 164175
rect -340 164147 -306 164175
rect -278 164147 -244 164175
rect -216 164147 -168 164175
rect -478 164113 -168 164147
rect -478 164085 -430 164113
rect -402 164085 -368 164113
rect -340 164085 -306 164113
rect -278 164085 -244 164113
rect -216 164085 -168 164113
rect -478 164051 -168 164085
rect -478 164023 -430 164051
rect -402 164023 -368 164051
rect -340 164023 -306 164051
rect -278 164023 -244 164051
rect -216 164023 -168 164051
rect -478 163989 -168 164023
rect -478 163961 -430 163989
rect -402 163961 -368 163989
rect -340 163961 -306 163989
rect -278 163961 -244 163989
rect -216 163961 -168 163989
rect -478 155175 -168 163961
rect 2086 286538 2114 286543
rect 2086 155554 2114 286510
rect 2709 281175 3019 289961
rect 2709 281147 2757 281175
rect 2785 281147 2819 281175
rect 2847 281147 2881 281175
rect 2909 281147 2943 281175
rect 2971 281147 3019 281175
rect 2709 281113 3019 281147
rect 2709 281085 2757 281113
rect 2785 281085 2819 281113
rect 2847 281085 2881 281113
rect 2909 281085 2943 281113
rect 2971 281085 3019 281113
rect 2709 281051 3019 281085
rect 2709 281023 2757 281051
rect 2785 281023 2819 281051
rect 2847 281023 2881 281051
rect 2909 281023 2943 281051
rect 2971 281023 3019 281051
rect 2709 280989 3019 281023
rect 2709 280961 2757 280989
rect 2785 280961 2819 280989
rect 2847 280961 2881 280989
rect 2909 280961 2943 280989
rect 2971 280961 3019 280989
rect 2709 272175 3019 280961
rect 3766 293594 3794 293599
rect 2709 272147 2757 272175
rect 2785 272147 2819 272175
rect 2847 272147 2881 272175
rect 2909 272147 2943 272175
rect 2971 272147 3019 272175
rect 2709 272113 3019 272147
rect 2709 272085 2757 272113
rect 2785 272085 2819 272113
rect 2847 272085 2881 272113
rect 2909 272085 2943 272113
rect 2971 272085 3019 272113
rect 2709 272051 3019 272085
rect 2709 272023 2757 272051
rect 2785 272023 2819 272051
rect 2847 272023 2881 272051
rect 2909 272023 2943 272051
rect 2971 272023 3019 272051
rect 2709 271989 3019 272023
rect 2709 271961 2757 271989
rect 2785 271961 2819 271989
rect 2847 271961 2881 271989
rect 2909 271961 2943 271989
rect 2971 271961 3019 271989
rect 2086 155521 2114 155526
rect 2142 265370 2170 265375
rect -478 155147 -430 155175
rect -402 155147 -368 155175
rect -340 155147 -306 155175
rect -278 155147 -244 155175
rect -216 155147 -168 155175
rect -478 155113 -168 155147
rect -478 155085 -430 155113
rect -402 155085 -368 155113
rect -340 155085 -306 155113
rect -278 155085 -244 155113
rect -216 155085 -168 155113
rect -478 155051 -168 155085
rect -478 155023 -430 155051
rect -402 155023 -368 155051
rect -340 155023 -306 155051
rect -278 155023 -244 155051
rect -216 155023 -168 155051
rect -478 154989 -168 155023
rect -478 154961 -430 154989
rect -402 154961 -368 154989
rect -340 154961 -306 154989
rect -278 154961 -244 154989
rect -216 154961 -168 154989
rect -478 146175 -168 154961
rect 2142 153874 2170 265342
rect 2709 263175 3019 271961
rect 2709 263147 2757 263175
rect 2785 263147 2819 263175
rect 2847 263147 2881 263175
rect 2909 263147 2943 263175
rect 2971 263147 3019 263175
rect 2709 263113 3019 263147
rect 2709 263085 2757 263113
rect 2785 263085 2819 263113
rect 2847 263085 2881 263113
rect 2909 263085 2943 263113
rect 2971 263085 3019 263113
rect 2709 263051 3019 263085
rect 2709 263023 2757 263051
rect 2785 263023 2819 263051
rect 2847 263023 2881 263051
rect 2909 263023 2943 263051
rect 2971 263023 3019 263051
rect 2709 262989 3019 263023
rect 2709 262961 2757 262989
rect 2785 262961 2819 262989
rect 2847 262961 2881 262989
rect 2909 262961 2943 262989
rect 2971 262961 3019 262989
rect 2709 254175 3019 262961
rect 2709 254147 2757 254175
rect 2785 254147 2819 254175
rect 2847 254147 2881 254175
rect 2909 254147 2943 254175
rect 2971 254147 3019 254175
rect 2709 254113 3019 254147
rect 2709 254085 2757 254113
rect 2785 254085 2819 254113
rect 2847 254085 2881 254113
rect 2909 254085 2943 254113
rect 2971 254085 3019 254113
rect 2709 254051 3019 254085
rect 2709 254023 2757 254051
rect 2785 254023 2819 254051
rect 2847 254023 2881 254051
rect 2909 254023 2943 254051
rect 2971 254023 3019 254051
rect 2709 253989 3019 254023
rect 2709 253961 2757 253989
rect 2785 253961 2819 253989
rect 2847 253961 2881 253989
rect 2909 253961 2943 253989
rect 2971 253961 3019 253989
rect 2709 245175 3019 253961
rect 2709 245147 2757 245175
rect 2785 245147 2819 245175
rect 2847 245147 2881 245175
rect 2909 245147 2943 245175
rect 2971 245147 3019 245175
rect 2709 245113 3019 245147
rect 2709 245085 2757 245113
rect 2785 245085 2819 245113
rect 2847 245085 2881 245113
rect 2909 245085 2943 245113
rect 2971 245085 3019 245113
rect 2709 245051 3019 245085
rect 2709 245023 2757 245051
rect 2785 245023 2819 245051
rect 2847 245023 2881 245051
rect 2909 245023 2943 245051
rect 2971 245023 3019 245051
rect 2709 244989 3019 245023
rect 2709 244961 2757 244989
rect 2785 244961 2819 244989
rect 2847 244961 2881 244989
rect 2909 244961 2943 244989
rect 2971 244961 3019 244989
rect 2142 153841 2170 153846
rect 2198 244202 2226 244207
rect -478 146147 -430 146175
rect -402 146147 -368 146175
rect -340 146147 -306 146175
rect -278 146147 -244 146175
rect -216 146147 -168 146175
rect -478 146113 -168 146147
rect -478 146085 -430 146113
rect -402 146085 -368 146113
rect -340 146085 -306 146113
rect -278 146085 -244 146113
rect -216 146085 -168 146113
rect -478 146051 -168 146085
rect -478 146023 -430 146051
rect -402 146023 -368 146051
rect -340 146023 -306 146051
rect -278 146023 -244 146051
rect -216 146023 -168 146051
rect -478 145989 -168 146023
rect -478 145961 -430 145989
rect -402 145961 -368 145989
rect -340 145961 -306 145989
rect -278 145961 -244 145989
rect -216 145961 -168 145989
rect -478 137175 -168 145961
rect 2086 152474 2114 152479
rect 2086 144914 2114 152446
rect 2198 152194 2226 244174
rect 2709 236175 3019 244961
rect 2709 236147 2757 236175
rect 2785 236147 2819 236175
rect 2847 236147 2881 236175
rect 2909 236147 2943 236175
rect 2971 236147 3019 236175
rect 2709 236113 3019 236147
rect 2709 236085 2757 236113
rect 2785 236085 2819 236113
rect 2847 236085 2881 236113
rect 2909 236085 2943 236113
rect 2971 236085 3019 236113
rect 2709 236051 3019 236085
rect 2709 236023 2757 236051
rect 2785 236023 2819 236051
rect 2847 236023 2881 236051
rect 2909 236023 2943 236051
rect 2971 236023 3019 236051
rect 2709 235989 3019 236023
rect 2709 235961 2757 235989
rect 2785 235961 2819 235989
rect 2847 235961 2881 235989
rect 2909 235961 2943 235989
rect 2971 235961 3019 235989
rect 2709 227175 3019 235961
rect 2709 227147 2757 227175
rect 2785 227147 2819 227175
rect 2847 227147 2881 227175
rect 2909 227147 2943 227175
rect 2971 227147 3019 227175
rect 2709 227113 3019 227147
rect 2709 227085 2757 227113
rect 2785 227085 2819 227113
rect 2847 227085 2881 227113
rect 2909 227085 2943 227113
rect 2971 227085 3019 227113
rect 2709 227051 3019 227085
rect 2709 227023 2757 227051
rect 2785 227023 2819 227051
rect 2847 227023 2881 227051
rect 2909 227023 2943 227051
rect 2971 227023 3019 227051
rect 2709 226989 3019 227023
rect 2709 226961 2757 226989
rect 2785 226961 2819 226989
rect 2847 226961 2881 226989
rect 2909 226961 2943 226989
rect 2971 226961 3019 226989
rect 2198 152161 2226 152166
rect 2254 223034 2282 223039
rect 2254 150514 2282 223006
rect 2709 218175 3019 226961
rect 2709 218147 2757 218175
rect 2785 218147 2819 218175
rect 2847 218147 2881 218175
rect 2909 218147 2943 218175
rect 2971 218147 3019 218175
rect 2709 218113 3019 218147
rect 2709 218085 2757 218113
rect 2785 218085 2819 218113
rect 2847 218085 2881 218113
rect 2909 218085 2943 218113
rect 2971 218085 3019 218113
rect 2709 218051 3019 218085
rect 2709 218023 2757 218051
rect 2785 218023 2819 218051
rect 2847 218023 2881 218051
rect 2909 218023 2943 218051
rect 2971 218023 3019 218051
rect 2709 217989 3019 218023
rect 2709 217961 2757 217989
rect 2785 217961 2819 217989
rect 2847 217961 2881 217989
rect 2909 217961 2943 217989
rect 2971 217961 3019 217989
rect 2709 209175 3019 217961
rect 2709 209147 2757 209175
rect 2785 209147 2819 209175
rect 2847 209147 2881 209175
rect 2909 209147 2943 209175
rect 2971 209147 3019 209175
rect 2709 209113 3019 209147
rect 2709 209085 2757 209113
rect 2785 209085 2819 209113
rect 2847 209085 2881 209113
rect 2909 209085 2943 209113
rect 2971 209085 3019 209113
rect 2709 209051 3019 209085
rect 2709 209023 2757 209051
rect 2785 209023 2819 209051
rect 2847 209023 2881 209051
rect 2909 209023 2943 209051
rect 2971 209023 3019 209051
rect 2709 208989 3019 209023
rect 2709 208961 2757 208989
rect 2785 208961 2819 208989
rect 2847 208961 2881 208989
rect 2909 208961 2943 208989
rect 2971 208961 3019 208989
rect 2709 200175 3019 208961
rect 2709 200147 2757 200175
rect 2785 200147 2819 200175
rect 2847 200147 2881 200175
rect 2909 200147 2943 200175
rect 2971 200147 3019 200175
rect 2709 200113 3019 200147
rect 2709 200085 2757 200113
rect 2785 200085 2819 200113
rect 2847 200085 2881 200113
rect 2909 200085 2943 200113
rect 2971 200085 3019 200113
rect 2709 200051 3019 200085
rect 2709 200023 2757 200051
rect 2785 200023 2819 200051
rect 2847 200023 2881 200051
rect 2909 200023 2943 200051
rect 2971 200023 3019 200051
rect 2709 199989 3019 200023
rect 2709 199961 2757 199989
rect 2785 199961 2819 199989
rect 2847 199961 2881 199989
rect 2909 199961 2943 199989
rect 2971 199961 3019 199989
rect 2709 191175 3019 199961
rect 2709 191147 2757 191175
rect 2785 191147 2819 191175
rect 2847 191147 2881 191175
rect 2909 191147 2943 191175
rect 2971 191147 3019 191175
rect 2709 191113 3019 191147
rect 2709 191085 2757 191113
rect 2785 191085 2819 191113
rect 2847 191085 2881 191113
rect 2909 191085 2943 191113
rect 2971 191085 3019 191113
rect 2709 191051 3019 191085
rect 2709 191023 2757 191051
rect 2785 191023 2819 191051
rect 2847 191023 2881 191051
rect 2909 191023 2943 191051
rect 2971 191023 3019 191051
rect 2709 190989 3019 191023
rect 2709 190961 2757 190989
rect 2785 190961 2819 190989
rect 2847 190961 2881 190989
rect 2909 190961 2943 190989
rect 2971 190961 3019 190989
rect 2709 182175 3019 190961
rect 2709 182147 2757 182175
rect 2785 182147 2819 182175
rect 2847 182147 2881 182175
rect 2909 182147 2943 182175
rect 2971 182147 3019 182175
rect 2709 182113 3019 182147
rect 2709 182085 2757 182113
rect 2785 182085 2819 182113
rect 2847 182085 2881 182113
rect 2909 182085 2943 182113
rect 2971 182085 3019 182113
rect 2709 182051 3019 182085
rect 2709 182023 2757 182051
rect 2785 182023 2819 182051
rect 2847 182023 2881 182051
rect 2909 182023 2943 182051
rect 2971 182023 3019 182051
rect 2709 181989 3019 182023
rect 2709 181961 2757 181989
rect 2785 181961 2819 181989
rect 2847 181961 2881 181989
rect 2909 181961 2943 181989
rect 2971 181961 3019 181989
rect 2254 150481 2282 150486
rect 2310 180698 2338 180703
rect 2310 147154 2338 180670
rect 2310 147121 2338 147126
rect 2709 173175 3019 181961
rect 2709 173147 2757 173175
rect 2785 173147 2819 173175
rect 2847 173147 2881 173175
rect 2909 173147 2943 173175
rect 2971 173147 3019 173175
rect 2709 173113 3019 173147
rect 2709 173085 2757 173113
rect 2785 173085 2819 173113
rect 2847 173085 2881 173113
rect 2909 173085 2943 173113
rect 2971 173085 3019 173113
rect 2709 173051 3019 173085
rect 2709 173023 2757 173051
rect 2785 173023 2819 173051
rect 2847 173023 2881 173051
rect 2909 173023 2943 173051
rect 2971 173023 3019 173051
rect 2709 172989 3019 173023
rect 2709 172961 2757 172989
rect 2785 172961 2819 172989
rect 2847 172961 2881 172989
rect 2909 172961 2943 172989
rect 2971 172961 3019 172989
rect 2709 164175 3019 172961
rect 2709 164147 2757 164175
rect 2785 164147 2819 164175
rect 2847 164147 2881 164175
rect 2909 164147 2943 164175
rect 2971 164147 3019 164175
rect 2709 164113 3019 164147
rect 2709 164085 2757 164113
rect 2785 164085 2819 164113
rect 2847 164085 2881 164113
rect 2909 164085 2943 164113
rect 2971 164085 3019 164113
rect 2709 164051 3019 164085
rect 2709 164023 2757 164051
rect 2785 164023 2819 164051
rect 2847 164023 2881 164051
rect 2909 164023 2943 164051
rect 2971 164023 3019 164051
rect 2709 163989 3019 164023
rect 2709 163961 2757 163989
rect 2785 163961 2819 163989
rect 2847 163961 2881 163989
rect 2909 163961 2943 163989
rect 2971 163961 3019 163989
rect 2709 155175 3019 163961
rect 2709 155147 2757 155175
rect 2785 155147 2819 155175
rect 2847 155147 2881 155175
rect 2909 155147 2943 155175
rect 2971 155147 3019 155175
rect 2709 155113 3019 155147
rect 2709 155085 2757 155113
rect 2785 155085 2819 155113
rect 2847 155085 2881 155113
rect 2909 155085 2943 155113
rect 2971 155085 3019 155113
rect 2709 155051 3019 155085
rect 2709 155023 2757 155051
rect 2785 155023 2819 155051
rect 2847 155023 2881 155051
rect 2909 155023 2943 155051
rect 2971 155023 3019 155051
rect 2709 154989 3019 155023
rect 2709 154961 2757 154989
rect 2785 154961 2819 154989
rect 2847 154961 2881 154989
rect 2909 154961 2943 154989
rect 2971 154961 3019 154989
rect 2709 146175 3019 154961
rect 3094 272426 3122 272431
rect 3094 154434 3122 272398
rect 3094 154401 3122 154406
rect 3150 173642 3178 173647
rect 3150 146594 3178 173614
rect 3766 156114 3794 293566
rect 4569 293175 4879 298872
rect 4569 293147 4617 293175
rect 4645 293147 4679 293175
rect 4707 293147 4741 293175
rect 4769 293147 4803 293175
rect 4831 293147 4879 293175
rect 4569 293113 4879 293147
rect 4569 293085 4617 293113
rect 4645 293085 4679 293113
rect 4707 293085 4741 293113
rect 4769 293085 4803 293113
rect 4831 293085 4879 293113
rect 4569 293051 4879 293085
rect 4569 293023 4617 293051
rect 4645 293023 4679 293051
rect 4707 293023 4741 293051
rect 4769 293023 4803 293051
rect 4831 293023 4879 293051
rect 4569 292989 4879 293023
rect 4569 292961 4617 292989
rect 4645 292961 4679 292989
rect 4707 292961 4741 292989
rect 4769 292961 4803 292989
rect 4831 292961 4879 292989
rect 4569 284175 4879 292961
rect 4569 284147 4617 284175
rect 4645 284147 4679 284175
rect 4707 284147 4741 284175
rect 4769 284147 4803 284175
rect 4831 284147 4879 284175
rect 4569 284113 4879 284147
rect 4569 284085 4617 284113
rect 4645 284085 4679 284113
rect 4707 284085 4741 284113
rect 4769 284085 4803 284113
rect 4831 284085 4879 284113
rect 4569 284051 4879 284085
rect 4569 284023 4617 284051
rect 4645 284023 4679 284051
rect 4707 284023 4741 284051
rect 4769 284023 4803 284051
rect 4831 284023 4879 284051
rect 4569 283989 4879 284023
rect 4569 283961 4617 283989
rect 4645 283961 4679 283989
rect 4707 283961 4741 283989
rect 4769 283961 4803 283989
rect 4831 283961 4879 283989
rect 4569 275175 4879 283961
rect 18069 298606 18379 299134
rect 18069 298578 18117 298606
rect 18145 298578 18179 298606
rect 18207 298578 18241 298606
rect 18269 298578 18303 298606
rect 18331 298578 18379 298606
rect 18069 298544 18379 298578
rect 18069 298516 18117 298544
rect 18145 298516 18179 298544
rect 18207 298516 18241 298544
rect 18269 298516 18303 298544
rect 18331 298516 18379 298544
rect 18069 298482 18379 298516
rect 18069 298454 18117 298482
rect 18145 298454 18179 298482
rect 18207 298454 18241 298482
rect 18269 298454 18303 298482
rect 18331 298454 18379 298482
rect 18069 298420 18379 298454
rect 18069 298392 18117 298420
rect 18145 298392 18179 298420
rect 18207 298392 18241 298420
rect 18269 298392 18303 298420
rect 18331 298392 18379 298420
rect 18069 290175 18379 298392
rect 18069 290147 18117 290175
rect 18145 290147 18179 290175
rect 18207 290147 18241 290175
rect 18269 290147 18303 290175
rect 18331 290147 18379 290175
rect 18069 290113 18379 290147
rect 18069 290085 18117 290113
rect 18145 290085 18179 290113
rect 18207 290085 18241 290113
rect 18269 290085 18303 290113
rect 18331 290085 18379 290113
rect 18069 290051 18379 290085
rect 18069 290023 18117 290051
rect 18145 290023 18179 290051
rect 18207 290023 18241 290051
rect 18269 290023 18303 290051
rect 18331 290023 18379 290051
rect 18069 289989 18379 290023
rect 18069 289961 18117 289989
rect 18145 289961 18179 289989
rect 18207 289961 18241 289989
rect 18269 289961 18303 289989
rect 18331 289961 18379 289989
rect 18069 281175 18379 289961
rect 18069 281147 18117 281175
rect 18145 281147 18179 281175
rect 18207 281147 18241 281175
rect 18269 281147 18303 281175
rect 18331 281147 18379 281175
rect 18069 281113 18379 281147
rect 18069 281085 18117 281113
rect 18145 281085 18179 281113
rect 18207 281085 18241 281113
rect 18269 281085 18303 281113
rect 18331 281085 18379 281113
rect 18069 281051 18379 281085
rect 18069 281023 18117 281051
rect 18145 281023 18179 281051
rect 18207 281023 18241 281051
rect 18269 281023 18303 281051
rect 18331 281023 18379 281051
rect 18069 280989 18379 281023
rect 18069 280961 18117 280989
rect 18145 280961 18179 280989
rect 18207 280961 18241 280989
rect 18269 280961 18303 280989
rect 18331 280961 18379 280989
rect 4569 275147 4617 275175
rect 4645 275147 4679 275175
rect 4707 275147 4741 275175
rect 4769 275147 4803 275175
rect 4831 275147 4879 275175
rect 4569 275113 4879 275147
rect 4569 275085 4617 275113
rect 4645 275085 4679 275113
rect 4707 275085 4741 275113
rect 4769 275085 4803 275113
rect 4831 275085 4879 275113
rect 4569 275051 4879 275085
rect 4569 275023 4617 275051
rect 4645 275023 4679 275051
rect 4707 275023 4741 275051
rect 4769 275023 4803 275051
rect 4831 275023 4879 275051
rect 4569 274989 4879 275023
rect 4569 274961 4617 274989
rect 4645 274961 4679 274989
rect 4707 274961 4741 274989
rect 4769 274961 4803 274989
rect 4831 274961 4879 274989
rect 4569 266175 4879 274961
rect 4569 266147 4617 266175
rect 4645 266147 4679 266175
rect 4707 266147 4741 266175
rect 4769 266147 4803 266175
rect 4831 266147 4879 266175
rect 4569 266113 4879 266147
rect 4569 266085 4617 266113
rect 4645 266085 4679 266113
rect 4707 266085 4741 266113
rect 4769 266085 4803 266113
rect 4831 266085 4879 266113
rect 4569 266051 4879 266085
rect 4569 266023 4617 266051
rect 4645 266023 4679 266051
rect 4707 266023 4741 266051
rect 4769 266023 4803 266051
rect 4831 266023 4879 266051
rect 4569 265989 4879 266023
rect 4569 265961 4617 265989
rect 4645 265961 4679 265989
rect 4707 265961 4741 265989
rect 4769 265961 4803 265989
rect 4831 265961 4879 265989
rect 4569 257175 4879 265961
rect 4569 257147 4617 257175
rect 4645 257147 4679 257175
rect 4707 257147 4741 257175
rect 4769 257147 4803 257175
rect 4831 257147 4879 257175
rect 4569 257113 4879 257147
rect 4569 257085 4617 257113
rect 4645 257085 4679 257113
rect 4707 257085 4741 257113
rect 4769 257085 4803 257113
rect 4831 257085 4879 257113
rect 4569 257051 4879 257085
rect 4569 257023 4617 257051
rect 4645 257023 4679 257051
rect 4707 257023 4741 257051
rect 4769 257023 4803 257051
rect 4831 257023 4879 257051
rect 4569 256989 4879 257023
rect 4569 256961 4617 256989
rect 4645 256961 4679 256989
rect 4707 256961 4741 256989
rect 4769 256961 4803 256989
rect 4831 256961 4879 256989
rect 3766 156081 3794 156086
rect 3822 251258 3850 251263
rect 3822 152754 3850 251230
rect 4569 248175 4879 256961
rect 4569 248147 4617 248175
rect 4645 248147 4679 248175
rect 4707 248147 4741 248175
rect 4769 248147 4803 248175
rect 4831 248147 4879 248175
rect 4569 248113 4879 248147
rect 4569 248085 4617 248113
rect 4645 248085 4679 248113
rect 4707 248085 4741 248113
rect 4769 248085 4803 248113
rect 4831 248085 4879 248113
rect 4569 248051 4879 248085
rect 4569 248023 4617 248051
rect 4645 248023 4679 248051
rect 4707 248023 4741 248051
rect 4769 248023 4803 248051
rect 4831 248023 4879 248051
rect 4569 247989 4879 248023
rect 4569 247961 4617 247989
rect 4645 247961 4679 247989
rect 4707 247961 4741 247989
rect 4769 247961 4803 247989
rect 4831 247961 4879 247989
rect 4569 239175 4879 247961
rect 4569 239147 4617 239175
rect 4645 239147 4679 239175
rect 4707 239147 4741 239175
rect 4769 239147 4803 239175
rect 4831 239147 4879 239175
rect 4569 239113 4879 239147
rect 4569 239085 4617 239113
rect 4645 239085 4679 239113
rect 4707 239085 4741 239113
rect 4769 239085 4803 239113
rect 4831 239085 4879 239113
rect 4569 239051 4879 239085
rect 4569 239023 4617 239051
rect 4645 239023 4679 239051
rect 4707 239023 4741 239051
rect 4769 239023 4803 239051
rect 4831 239023 4879 239051
rect 4569 238989 4879 239023
rect 4569 238961 4617 238989
rect 4645 238961 4679 238989
rect 4707 238961 4741 238989
rect 4769 238961 4803 238989
rect 4831 238961 4879 238989
rect 4569 230175 4879 238961
rect 4569 230147 4617 230175
rect 4645 230147 4679 230175
rect 4707 230147 4741 230175
rect 4769 230147 4803 230175
rect 4831 230147 4879 230175
rect 4569 230113 4879 230147
rect 3822 152721 3850 152726
rect 3878 230090 3906 230095
rect 3878 151074 3906 230062
rect 4569 230085 4617 230113
rect 4645 230085 4679 230113
rect 4707 230085 4741 230113
rect 4769 230085 4803 230113
rect 4831 230085 4879 230113
rect 4569 230051 4879 230085
rect 4569 230023 4617 230051
rect 4645 230023 4679 230051
rect 4707 230023 4741 230051
rect 4769 230023 4803 230051
rect 4831 230023 4879 230051
rect 4569 229989 4879 230023
rect 4569 229961 4617 229989
rect 4645 229961 4679 229989
rect 4707 229961 4741 229989
rect 4769 229961 4803 229989
rect 4831 229961 4879 229989
rect 4569 221175 4879 229961
rect 4569 221147 4617 221175
rect 4645 221147 4679 221175
rect 4707 221147 4741 221175
rect 4769 221147 4803 221175
rect 4831 221147 4879 221175
rect 4569 221113 4879 221147
rect 4569 221085 4617 221113
rect 4645 221085 4679 221113
rect 4707 221085 4741 221113
rect 4769 221085 4803 221113
rect 4831 221085 4879 221113
rect 4569 221051 4879 221085
rect 4569 221023 4617 221051
rect 4645 221023 4679 221051
rect 4707 221023 4741 221051
rect 4769 221023 4803 221051
rect 4831 221023 4879 221051
rect 4569 220989 4879 221023
rect 4569 220961 4617 220989
rect 4645 220961 4679 220989
rect 4707 220961 4741 220989
rect 4769 220961 4803 220989
rect 4831 220961 4879 220989
rect 4569 212175 4879 220961
rect 4569 212147 4617 212175
rect 4645 212147 4679 212175
rect 4707 212147 4741 212175
rect 4769 212147 4803 212175
rect 4831 212147 4879 212175
rect 4569 212113 4879 212147
rect 4569 212085 4617 212113
rect 4645 212085 4679 212113
rect 4707 212085 4741 212113
rect 4769 212085 4803 212113
rect 4831 212085 4879 212113
rect 4569 212051 4879 212085
rect 4569 212023 4617 212051
rect 4645 212023 4679 212051
rect 4707 212023 4741 212051
rect 4769 212023 4803 212051
rect 4831 212023 4879 212051
rect 4569 211989 4879 212023
rect 4569 211961 4617 211989
rect 4645 211961 4679 211989
rect 4707 211961 4741 211989
rect 4769 211961 4803 211989
rect 4831 211961 4879 211989
rect 3878 151041 3906 151046
rect 3934 208922 3962 208927
rect 3934 149394 3962 208894
rect 4569 203175 4879 211961
rect 4569 203147 4617 203175
rect 4645 203147 4679 203175
rect 4707 203147 4741 203175
rect 4769 203147 4803 203175
rect 4831 203147 4879 203175
rect 4569 203113 4879 203147
rect 4569 203085 4617 203113
rect 4645 203085 4679 203113
rect 4707 203085 4741 203113
rect 4769 203085 4803 203113
rect 4831 203085 4879 203113
rect 4569 203051 4879 203085
rect 4569 203023 4617 203051
rect 4645 203023 4679 203051
rect 4707 203023 4741 203051
rect 4769 203023 4803 203051
rect 4831 203023 4879 203051
rect 4569 202989 4879 203023
rect 4569 202961 4617 202989
rect 4645 202961 4679 202989
rect 4707 202961 4741 202989
rect 4769 202961 4803 202989
rect 4831 202961 4879 202989
rect 4569 194175 4879 202961
rect 4569 194147 4617 194175
rect 4645 194147 4679 194175
rect 4707 194147 4741 194175
rect 4769 194147 4803 194175
rect 4831 194147 4879 194175
rect 4569 194113 4879 194147
rect 4569 194085 4617 194113
rect 4645 194085 4679 194113
rect 4707 194085 4741 194113
rect 4769 194085 4803 194113
rect 4831 194085 4879 194113
rect 4569 194051 4879 194085
rect 4569 194023 4617 194051
rect 4645 194023 4679 194051
rect 4707 194023 4741 194051
rect 4769 194023 4803 194051
rect 4831 194023 4879 194051
rect 4569 193989 4879 194023
rect 4569 193961 4617 193989
rect 4645 193961 4679 193989
rect 4707 193961 4741 193989
rect 4769 193961 4803 193989
rect 4831 193961 4879 193989
rect 4569 185175 4879 193961
rect 5446 279482 5474 279487
rect 4569 185147 4617 185175
rect 4645 185147 4679 185175
rect 4707 185147 4741 185175
rect 4769 185147 4803 185175
rect 4831 185147 4879 185175
rect 4569 185113 4879 185147
rect 4569 185085 4617 185113
rect 4645 185085 4679 185113
rect 4707 185085 4741 185113
rect 4769 185085 4803 185113
rect 4831 185085 4879 185113
rect 4569 185051 4879 185085
rect 4569 185023 4617 185051
rect 4645 185023 4679 185051
rect 4707 185023 4741 185051
rect 4769 185023 4803 185051
rect 4831 185023 4879 185051
rect 4569 184989 4879 185023
rect 4569 184961 4617 184989
rect 4645 184961 4679 184989
rect 4707 184961 4741 184989
rect 4769 184961 4803 184989
rect 4831 184961 4879 184989
rect 4569 176175 4879 184961
rect 4569 176147 4617 176175
rect 4645 176147 4679 176175
rect 4707 176147 4741 176175
rect 4769 176147 4803 176175
rect 4831 176147 4879 176175
rect 4569 176113 4879 176147
rect 4569 176085 4617 176113
rect 4645 176085 4679 176113
rect 4707 176085 4741 176113
rect 4769 176085 4803 176113
rect 4831 176085 4879 176113
rect 4569 176051 4879 176085
rect 4569 176023 4617 176051
rect 4645 176023 4679 176051
rect 4707 176023 4741 176051
rect 4769 176023 4803 176051
rect 4831 176023 4879 176051
rect 4569 175989 4879 176023
rect 4569 175961 4617 175989
rect 4645 175961 4679 175989
rect 4707 175961 4741 175989
rect 4769 175961 4803 175989
rect 4831 175961 4879 175989
rect 4569 167175 4879 175961
rect 4569 167147 4617 167175
rect 4645 167147 4679 167175
rect 4707 167147 4741 167175
rect 4769 167147 4803 167175
rect 4831 167147 4879 167175
rect 4569 167113 4879 167147
rect 4569 167085 4617 167113
rect 4645 167085 4679 167113
rect 4707 167085 4741 167113
rect 4769 167085 4803 167113
rect 4831 167085 4879 167113
rect 4569 167051 4879 167085
rect 4569 167023 4617 167051
rect 4645 167023 4679 167051
rect 4707 167023 4741 167051
rect 4769 167023 4803 167051
rect 4831 167023 4879 167051
rect 4569 166989 4879 167023
rect 4569 166961 4617 166989
rect 4645 166961 4679 166989
rect 4707 166961 4741 166989
rect 4769 166961 4803 166989
rect 4831 166961 4879 166989
rect 3934 149361 3962 149366
rect 3990 166586 4018 166591
rect 3150 146561 3178 146566
rect 2709 146147 2757 146175
rect 2785 146147 2819 146175
rect 2847 146147 2881 146175
rect 2909 146147 2943 146175
rect 2971 146147 3019 146175
rect 2709 146113 3019 146147
rect 2709 146085 2757 146113
rect 2785 146085 2819 146113
rect 2847 146085 2881 146113
rect 2909 146085 2943 146113
rect 2971 146085 3019 146113
rect 2709 146051 3019 146085
rect 2709 146023 2757 146051
rect 2785 146023 2819 146051
rect 2847 146023 2881 146051
rect 2909 146023 2943 146051
rect 2971 146023 3019 146051
rect 2709 145989 3019 146023
rect 3990 146034 4018 166558
rect 3990 146001 4018 146006
rect 4569 158175 4879 166961
rect 4569 158147 4617 158175
rect 4645 158147 4679 158175
rect 4707 158147 4741 158175
rect 4769 158147 4803 158175
rect 4831 158147 4879 158175
rect 4569 158113 4879 158147
rect 4569 158085 4617 158113
rect 4645 158085 4679 158113
rect 4707 158085 4741 158113
rect 4769 158085 4803 158113
rect 4831 158085 4879 158113
rect 4569 158051 4879 158085
rect 4569 158023 4617 158051
rect 4645 158023 4679 158051
rect 4707 158023 4741 158051
rect 4769 158023 4803 158051
rect 4831 158023 4879 158051
rect 4569 157989 4879 158023
rect 4569 157961 4617 157989
rect 4645 157961 4679 157989
rect 4707 157961 4741 157989
rect 4769 157961 4803 157989
rect 4831 157961 4879 157989
rect 4569 149175 4879 157961
rect 4569 149147 4617 149175
rect 4645 149147 4679 149175
rect 4707 149147 4741 149175
rect 4769 149147 4803 149175
rect 4831 149147 4879 149175
rect 4569 149113 4879 149147
rect 4569 149085 4617 149113
rect 4645 149085 4679 149113
rect 4707 149085 4741 149113
rect 4769 149085 4803 149113
rect 4831 149085 4879 149113
rect 4569 149051 4879 149085
rect 4569 149023 4617 149051
rect 4645 149023 4679 149051
rect 4707 149023 4741 149051
rect 4769 149023 4803 149051
rect 4831 149023 4879 149051
rect 4569 148989 4879 149023
rect 4569 148961 4617 148989
rect 4645 148961 4679 148989
rect 4707 148961 4741 148989
rect 4769 148961 4803 148989
rect 4831 148961 4879 148989
rect 2709 145961 2757 145989
rect 2785 145961 2819 145989
rect 2847 145961 2881 145989
rect 2909 145961 2943 145989
rect 2971 145961 3019 145989
rect 2086 144881 2114 144886
rect 2478 145418 2506 145423
rect 2478 144354 2506 145390
rect 2478 144321 2506 144326
rect 2086 143794 2114 143799
rect 2086 138474 2114 143766
rect 2086 138441 2114 138446
rect 2366 142114 2394 142119
rect -478 137147 -430 137175
rect -402 137147 -368 137175
rect -340 137147 -306 137175
rect -278 137147 -244 137175
rect -216 137147 -168 137175
rect -478 137113 -168 137147
rect -478 137085 -430 137113
rect -402 137085 -368 137113
rect -340 137085 -306 137113
rect -278 137085 -244 137113
rect -216 137085 -168 137113
rect -478 137051 -168 137085
rect 2310 138194 2338 138199
rect -478 137023 -430 137051
rect -402 137023 -368 137051
rect -340 137023 -306 137051
rect -278 137023 -244 137051
rect -216 137023 -168 137051
rect -478 136989 -168 137023
rect -478 136961 -430 136989
rect -402 136961 -368 136989
rect -340 136961 -306 136989
rect -278 136961 -244 136989
rect -216 136961 -168 136989
rect -478 128175 -168 136961
rect 2254 137074 2282 137079
rect 2198 136514 2226 136519
rect 2142 133714 2170 133719
rect -478 128147 -430 128175
rect -402 128147 -368 128175
rect -340 128147 -306 128175
rect -278 128147 -244 128175
rect -216 128147 -168 128175
rect -478 128113 -168 128147
rect -478 128085 -430 128113
rect -402 128085 -368 128113
rect -340 128085 -306 128113
rect -278 128085 -244 128113
rect -216 128085 -168 128113
rect -478 128051 -168 128085
rect -478 128023 -430 128051
rect -402 128023 -368 128051
rect -340 128023 -306 128051
rect -278 128023 -244 128051
rect -216 128023 -168 128051
rect -478 127989 -168 128023
rect -478 127961 -430 127989
rect -402 127961 -368 127989
rect -340 127961 -306 127989
rect -278 127961 -244 127989
rect -216 127961 -168 127989
rect -478 119175 -168 127961
rect -478 119147 -430 119175
rect -402 119147 -368 119175
rect -340 119147 -306 119175
rect -278 119147 -244 119175
rect -216 119147 -168 119175
rect -478 119113 -168 119147
rect -478 119085 -430 119113
rect -402 119085 -368 119113
rect -340 119085 -306 119113
rect -278 119085 -244 119113
rect -216 119085 -168 119113
rect -478 119051 -168 119085
rect -478 119023 -430 119051
rect -402 119023 -368 119051
rect -340 119023 -306 119051
rect -278 119023 -244 119051
rect -216 119023 -168 119051
rect -478 118989 -168 119023
rect -478 118961 -430 118989
rect -402 118961 -368 118989
rect -340 118961 -306 118989
rect -278 118961 -244 118989
rect -216 118961 -168 118989
rect -478 110175 -168 118961
rect -478 110147 -430 110175
rect -402 110147 -368 110175
rect -340 110147 -306 110175
rect -278 110147 -244 110175
rect -216 110147 -168 110175
rect -478 110113 -168 110147
rect -478 110085 -430 110113
rect -402 110085 -368 110113
rect -340 110085 -306 110113
rect -278 110085 -244 110113
rect -216 110085 -168 110113
rect -478 110051 -168 110085
rect -478 110023 -430 110051
rect -402 110023 -368 110051
rect -340 110023 -306 110051
rect -278 110023 -244 110051
rect -216 110023 -168 110051
rect -478 109989 -168 110023
rect -478 109961 -430 109989
rect -402 109961 -368 109989
rect -340 109961 -306 109989
rect -278 109961 -244 109989
rect -216 109961 -168 109989
rect -478 101175 -168 109961
rect -478 101147 -430 101175
rect -402 101147 -368 101175
rect -340 101147 -306 101175
rect -278 101147 -244 101175
rect -216 101147 -168 101175
rect -478 101113 -168 101147
rect -478 101085 -430 101113
rect -402 101085 -368 101113
rect -340 101085 -306 101113
rect -278 101085 -244 101113
rect -216 101085 -168 101113
rect -478 101051 -168 101085
rect -478 101023 -430 101051
rect -402 101023 -368 101051
rect -340 101023 -306 101051
rect -278 101023 -244 101051
rect -216 101023 -168 101051
rect -478 100989 -168 101023
rect -478 100961 -430 100989
rect -402 100961 -368 100989
rect -340 100961 -306 100989
rect -278 100961 -244 100989
rect -216 100961 -168 100989
rect -478 92175 -168 100961
rect -478 92147 -430 92175
rect -402 92147 -368 92175
rect -340 92147 -306 92175
rect -278 92147 -244 92175
rect -216 92147 -168 92175
rect -478 92113 -168 92147
rect -478 92085 -430 92113
rect -402 92085 -368 92113
rect -340 92085 -306 92113
rect -278 92085 -244 92113
rect -216 92085 -168 92113
rect -478 92051 -168 92085
rect -478 92023 -430 92051
rect -402 92023 -368 92051
rect -340 92023 -306 92051
rect -278 92023 -244 92051
rect -216 92023 -168 92051
rect -478 91989 -168 92023
rect -478 91961 -430 91989
rect -402 91961 -368 91989
rect -340 91961 -306 91989
rect -278 91961 -244 91989
rect -216 91961 -168 91989
rect -478 83175 -168 91961
rect -478 83147 -430 83175
rect -402 83147 -368 83175
rect -340 83147 -306 83175
rect -278 83147 -244 83175
rect -216 83147 -168 83175
rect -478 83113 -168 83147
rect -478 83085 -430 83113
rect -402 83085 -368 83113
rect -340 83085 -306 83113
rect -278 83085 -244 83113
rect -216 83085 -168 83113
rect -478 83051 -168 83085
rect -478 83023 -430 83051
rect -402 83023 -368 83051
rect -340 83023 -306 83051
rect -278 83023 -244 83051
rect -216 83023 -168 83051
rect -478 82989 -168 83023
rect -478 82961 -430 82989
rect -402 82961 -368 82989
rect -340 82961 -306 82989
rect -278 82961 -244 82989
rect -216 82961 -168 82989
rect -478 74175 -168 82961
rect -478 74147 -430 74175
rect -402 74147 -368 74175
rect -340 74147 -306 74175
rect -278 74147 -244 74175
rect -216 74147 -168 74175
rect -478 74113 -168 74147
rect -478 74085 -430 74113
rect -402 74085 -368 74113
rect -340 74085 -306 74113
rect -278 74085 -244 74113
rect -216 74085 -168 74113
rect -478 74051 -168 74085
rect -478 74023 -430 74051
rect -402 74023 -368 74051
rect -340 74023 -306 74051
rect -278 74023 -244 74051
rect -216 74023 -168 74051
rect -478 73989 -168 74023
rect -478 73961 -430 73989
rect -402 73961 -368 73989
rect -340 73961 -306 73989
rect -278 73961 -244 73989
rect -216 73961 -168 73989
rect -478 65175 -168 73961
rect -478 65147 -430 65175
rect -402 65147 -368 65175
rect -340 65147 -306 65175
rect -278 65147 -244 65175
rect -216 65147 -168 65175
rect -478 65113 -168 65147
rect -478 65085 -430 65113
rect -402 65085 -368 65113
rect -340 65085 -306 65113
rect -278 65085 -244 65113
rect -216 65085 -168 65113
rect -478 65051 -168 65085
rect -478 65023 -430 65051
rect -402 65023 -368 65051
rect -340 65023 -306 65051
rect -278 65023 -244 65051
rect -216 65023 -168 65051
rect -478 64989 -168 65023
rect -478 64961 -430 64989
rect -402 64961 -368 64989
rect -340 64961 -306 64989
rect -278 64961 -244 64989
rect -216 64961 -168 64989
rect -478 56175 -168 64961
rect -478 56147 -430 56175
rect -402 56147 -368 56175
rect -340 56147 -306 56175
rect -278 56147 -244 56175
rect -216 56147 -168 56175
rect -478 56113 -168 56147
rect -478 56085 -430 56113
rect -402 56085 -368 56113
rect -340 56085 -306 56113
rect -278 56085 -244 56113
rect -216 56085 -168 56113
rect -478 56051 -168 56085
rect -478 56023 -430 56051
rect -402 56023 -368 56051
rect -340 56023 -306 56051
rect -278 56023 -244 56051
rect -216 56023 -168 56051
rect -478 55989 -168 56023
rect -478 55961 -430 55989
rect -402 55961 -368 55989
rect -340 55961 -306 55989
rect -278 55961 -244 55989
rect -216 55961 -168 55989
rect -478 47175 -168 55961
rect -478 47147 -430 47175
rect -402 47147 -368 47175
rect -340 47147 -306 47175
rect -278 47147 -244 47175
rect -216 47147 -168 47175
rect -478 47113 -168 47147
rect -478 47085 -430 47113
rect -402 47085 -368 47113
rect -340 47085 -306 47113
rect -278 47085 -244 47113
rect -216 47085 -168 47113
rect -478 47051 -168 47085
rect -478 47023 -430 47051
rect -402 47023 -368 47051
rect -340 47023 -306 47051
rect -278 47023 -244 47051
rect -216 47023 -168 47051
rect -478 46989 -168 47023
rect -478 46961 -430 46989
rect -402 46961 -368 46989
rect -340 46961 -306 46989
rect -278 46961 -244 46989
rect -216 46961 -168 46989
rect -478 38175 -168 46961
rect -478 38147 -430 38175
rect -402 38147 -368 38175
rect -340 38147 -306 38175
rect -278 38147 -244 38175
rect -216 38147 -168 38175
rect -478 38113 -168 38147
rect -478 38085 -430 38113
rect -402 38085 -368 38113
rect -340 38085 -306 38113
rect -278 38085 -244 38113
rect -216 38085 -168 38113
rect -478 38051 -168 38085
rect -478 38023 -430 38051
rect -402 38023 -368 38051
rect -340 38023 -306 38051
rect -278 38023 -244 38051
rect -216 38023 -168 38051
rect -478 37989 -168 38023
rect -478 37961 -430 37989
rect -402 37961 -368 37989
rect -340 37961 -306 37989
rect -278 37961 -244 37989
rect -216 37961 -168 37989
rect -478 29175 -168 37961
rect -478 29147 -430 29175
rect -402 29147 -368 29175
rect -340 29147 -306 29175
rect -278 29147 -244 29175
rect -216 29147 -168 29175
rect -478 29113 -168 29147
rect -478 29085 -430 29113
rect -402 29085 -368 29113
rect -340 29085 -306 29113
rect -278 29085 -244 29113
rect -216 29085 -168 29113
rect -478 29051 -168 29085
rect -478 29023 -430 29051
rect -402 29023 -368 29051
rect -340 29023 -306 29051
rect -278 29023 -244 29051
rect -216 29023 -168 29051
rect -478 28989 -168 29023
rect -478 28961 -430 28989
rect -402 28961 -368 28989
rect -340 28961 -306 28989
rect -278 28961 -244 28989
rect -216 28961 -168 28989
rect -478 20175 -168 28961
rect -478 20147 -430 20175
rect -402 20147 -368 20175
rect -340 20147 -306 20175
rect -278 20147 -244 20175
rect -216 20147 -168 20175
rect -478 20113 -168 20147
rect -478 20085 -430 20113
rect -402 20085 -368 20113
rect -340 20085 -306 20113
rect -278 20085 -244 20113
rect -216 20085 -168 20113
rect -478 20051 -168 20085
rect -478 20023 -430 20051
rect -402 20023 -368 20051
rect -340 20023 -306 20051
rect -278 20023 -244 20051
rect -216 20023 -168 20051
rect -478 19989 -168 20023
rect -478 19961 -430 19989
rect -402 19961 -368 19989
rect -340 19961 -306 19989
rect -278 19961 -244 19989
rect -216 19961 -168 19989
rect -478 11175 -168 19961
rect -478 11147 -430 11175
rect -402 11147 -368 11175
rect -340 11147 -306 11175
rect -278 11147 -244 11175
rect -216 11147 -168 11175
rect -478 11113 -168 11147
rect -478 11085 -430 11113
rect -402 11085 -368 11113
rect -340 11085 -306 11113
rect -278 11085 -244 11113
rect -216 11085 -168 11113
rect -478 11051 -168 11085
rect -478 11023 -430 11051
rect -402 11023 -368 11051
rect -340 11023 -306 11051
rect -278 11023 -244 11051
rect -216 11023 -168 11051
rect -478 10989 -168 11023
rect -478 10961 -430 10989
rect -402 10961 -368 10989
rect -340 10961 -306 10989
rect -278 10961 -244 10989
rect -216 10961 -168 10989
rect -478 2175 -168 10961
rect 2086 133154 2114 133159
rect 2086 4410 2114 133126
rect 2142 11466 2170 133686
rect 2198 46746 2226 136486
rect 2254 53746 2282 137046
rect 2310 67914 2338 138166
rect 2366 117306 2394 142086
rect 2366 117273 2394 117278
rect 2709 137175 3019 145961
rect 2709 137147 2757 137175
rect 2785 137147 2819 137175
rect 2847 137147 2881 137175
rect 2909 137147 2943 137175
rect 2971 137147 3019 137175
rect 2709 137113 3019 137147
rect 2709 137085 2757 137113
rect 2785 137085 2819 137113
rect 2847 137085 2881 137113
rect 2909 137085 2943 137113
rect 2971 137085 3019 137113
rect 2709 137051 3019 137085
rect 2709 137023 2757 137051
rect 2785 137023 2819 137051
rect 2847 137023 2881 137051
rect 2909 137023 2943 137051
rect 2971 137023 3019 137051
rect 2709 136989 3019 137023
rect 2709 136961 2757 136989
rect 2785 136961 2819 136989
rect 2847 136961 2881 136989
rect 2909 136961 2943 136989
rect 2971 136961 3019 136989
rect 2709 128175 3019 136961
rect 3150 140994 3178 140999
rect 2709 128147 2757 128175
rect 2785 128147 2819 128175
rect 2847 128147 2881 128175
rect 2909 128147 2943 128175
rect 2971 128147 3019 128175
rect 2709 128113 3019 128147
rect 2709 128085 2757 128113
rect 2785 128085 2819 128113
rect 2847 128085 2881 128113
rect 2909 128085 2943 128113
rect 2971 128085 3019 128113
rect 2709 128051 3019 128085
rect 2709 128023 2757 128051
rect 2785 128023 2819 128051
rect 2847 128023 2881 128051
rect 2909 128023 2943 128051
rect 2971 128023 3019 128051
rect 2709 127989 3019 128023
rect 2709 127961 2757 127989
rect 2785 127961 2819 127989
rect 2847 127961 2881 127989
rect 2909 127961 2943 127989
rect 2971 127961 3019 127989
rect 2709 119175 3019 127961
rect 2709 119147 2757 119175
rect 2785 119147 2819 119175
rect 2847 119147 2881 119175
rect 2909 119147 2943 119175
rect 2971 119147 3019 119175
rect 2709 119113 3019 119147
rect 2709 119085 2757 119113
rect 2785 119085 2819 119113
rect 2847 119085 2881 119113
rect 2909 119085 2943 119113
rect 2971 119085 3019 119113
rect 2709 119051 3019 119085
rect 2709 119023 2757 119051
rect 2785 119023 2819 119051
rect 2847 119023 2881 119051
rect 2909 119023 2943 119051
rect 2971 119023 3019 119051
rect 2709 118989 3019 119023
rect 2709 118961 2757 118989
rect 2785 118961 2819 118989
rect 2847 118961 2881 118989
rect 2909 118961 2943 118989
rect 2971 118961 3019 118989
rect 2310 67881 2338 67886
rect 2709 110175 3019 118961
rect 2709 110147 2757 110175
rect 2785 110147 2819 110175
rect 2847 110147 2881 110175
rect 2909 110147 2943 110175
rect 2971 110147 3019 110175
rect 2709 110113 3019 110147
rect 2709 110085 2757 110113
rect 2785 110085 2819 110113
rect 2847 110085 2881 110113
rect 2909 110085 2943 110113
rect 2971 110085 3019 110113
rect 2709 110051 3019 110085
rect 2709 110023 2757 110051
rect 2785 110023 2819 110051
rect 2847 110023 2881 110051
rect 2909 110023 2943 110051
rect 2971 110023 3019 110051
rect 2709 109989 3019 110023
rect 2709 109961 2757 109989
rect 2785 109961 2819 109989
rect 2847 109961 2881 109989
rect 2909 109961 2943 109989
rect 2971 109961 3019 109989
rect 2709 101175 3019 109961
rect 2709 101147 2757 101175
rect 2785 101147 2819 101175
rect 2847 101147 2881 101175
rect 2909 101147 2943 101175
rect 2971 101147 3019 101175
rect 2709 101113 3019 101147
rect 2709 101085 2757 101113
rect 2785 101085 2819 101113
rect 2847 101085 2881 101113
rect 2909 101085 2943 101113
rect 2971 101085 3019 101113
rect 2709 101051 3019 101085
rect 2709 101023 2757 101051
rect 2785 101023 2819 101051
rect 2847 101023 2881 101051
rect 2909 101023 2943 101051
rect 2971 101023 3019 101051
rect 2709 100989 3019 101023
rect 2709 100961 2757 100989
rect 2785 100961 2819 100989
rect 2847 100961 2881 100989
rect 2909 100961 2943 100989
rect 2971 100961 3019 100989
rect 2709 92175 3019 100961
rect 2709 92147 2757 92175
rect 2785 92147 2819 92175
rect 2847 92147 2881 92175
rect 2909 92147 2943 92175
rect 2971 92147 3019 92175
rect 2709 92113 3019 92147
rect 2709 92085 2757 92113
rect 2785 92085 2819 92113
rect 2847 92085 2881 92113
rect 2909 92085 2943 92113
rect 2971 92085 3019 92113
rect 2709 92051 3019 92085
rect 2709 92023 2757 92051
rect 2785 92023 2819 92051
rect 2847 92023 2881 92051
rect 2909 92023 2943 92051
rect 2971 92023 3019 92051
rect 2709 91989 3019 92023
rect 2709 91961 2757 91989
rect 2785 91961 2819 91989
rect 2847 91961 2881 91989
rect 2909 91961 2943 91989
rect 2971 91961 3019 91989
rect 2709 83175 3019 91961
rect 2709 83147 2757 83175
rect 2785 83147 2819 83175
rect 2847 83147 2881 83175
rect 2909 83147 2943 83175
rect 2971 83147 3019 83175
rect 2709 83113 3019 83147
rect 2709 83085 2757 83113
rect 2785 83085 2819 83113
rect 2847 83085 2881 83113
rect 2909 83085 2943 83113
rect 2971 83085 3019 83113
rect 2709 83051 3019 83085
rect 2709 83023 2757 83051
rect 2785 83023 2819 83051
rect 2847 83023 2881 83051
rect 2909 83023 2943 83051
rect 2971 83023 3019 83051
rect 2709 82989 3019 83023
rect 2709 82961 2757 82989
rect 2785 82961 2819 82989
rect 2847 82961 2881 82989
rect 2909 82961 2943 82989
rect 2971 82961 3019 82989
rect 2709 74175 3019 82961
rect 2709 74147 2757 74175
rect 2785 74147 2819 74175
rect 2847 74147 2881 74175
rect 2909 74147 2943 74175
rect 2971 74147 3019 74175
rect 2709 74113 3019 74147
rect 2709 74085 2757 74113
rect 2785 74085 2819 74113
rect 2847 74085 2881 74113
rect 2909 74085 2943 74113
rect 2971 74085 3019 74113
rect 2709 74051 3019 74085
rect 2709 74023 2757 74051
rect 2785 74023 2819 74051
rect 2847 74023 2881 74051
rect 2909 74023 2943 74051
rect 2971 74023 3019 74051
rect 2709 73989 3019 74023
rect 2709 73961 2757 73989
rect 2785 73961 2819 73989
rect 2847 73961 2881 73989
rect 2909 73961 2943 73989
rect 2971 73961 3019 73989
rect 2254 53713 2282 53718
rect 2709 65175 3019 73961
rect 2709 65147 2757 65175
rect 2785 65147 2819 65175
rect 2847 65147 2881 65175
rect 2909 65147 2943 65175
rect 2971 65147 3019 65175
rect 2709 65113 3019 65147
rect 2709 65085 2757 65113
rect 2785 65085 2819 65113
rect 2847 65085 2881 65113
rect 2909 65085 2943 65113
rect 2971 65085 3019 65113
rect 2709 65051 3019 65085
rect 2709 65023 2757 65051
rect 2785 65023 2819 65051
rect 2847 65023 2881 65051
rect 2909 65023 2943 65051
rect 2971 65023 3019 65051
rect 2709 64989 3019 65023
rect 2709 64961 2757 64989
rect 2785 64961 2819 64989
rect 2847 64961 2881 64989
rect 2909 64961 2943 64989
rect 2971 64961 3019 64989
rect 2709 56175 3019 64961
rect 2709 56147 2757 56175
rect 2785 56147 2819 56175
rect 2847 56147 2881 56175
rect 2909 56147 2943 56175
rect 2971 56147 3019 56175
rect 2709 56113 3019 56147
rect 2709 56085 2757 56113
rect 2785 56085 2819 56113
rect 2847 56085 2881 56113
rect 2909 56085 2943 56113
rect 2971 56085 3019 56113
rect 2709 56051 3019 56085
rect 2709 56023 2757 56051
rect 2785 56023 2819 56051
rect 2847 56023 2881 56051
rect 2909 56023 2943 56051
rect 2971 56023 3019 56051
rect 2709 55989 3019 56023
rect 2709 55961 2757 55989
rect 2785 55961 2819 55989
rect 2847 55961 2881 55989
rect 2909 55961 2943 55989
rect 2971 55961 3019 55989
rect 2198 46713 2226 46718
rect 2709 47175 3019 55961
rect 2709 47147 2757 47175
rect 2785 47147 2819 47175
rect 2847 47147 2881 47175
rect 2909 47147 2943 47175
rect 2971 47147 3019 47175
rect 2709 47113 3019 47147
rect 2709 47085 2757 47113
rect 2785 47085 2819 47113
rect 2847 47085 2881 47113
rect 2909 47085 2943 47113
rect 2971 47085 3019 47113
rect 2709 47051 3019 47085
rect 2709 47023 2757 47051
rect 2785 47023 2819 47051
rect 2847 47023 2881 47051
rect 2909 47023 2943 47051
rect 2971 47023 3019 47051
rect 2709 46989 3019 47023
rect 2709 46961 2757 46989
rect 2785 46961 2819 46989
rect 2847 46961 2881 46989
rect 2909 46961 2943 46989
rect 2971 46961 3019 46989
rect 2142 11433 2170 11438
rect 2709 38175 3019 46961
rect 3094 135954 3122 135959
rect 3094 39690 3122 135926
rect 3150 103194 3178 140966
rect 4569 140175 4879 148961
rect 4942 187754 4970 187759
rect 4942 147714 4970 187726
rect 5446 154994 5474 279454
rect 18069 272175 18379 280961
rect 18069 272147 18117 272175
rect 18145 272147 18179 272175
rect 18207 272147 18241 272175
rect 18269 272147 18303 272175
rect 18331 272147 18379 272175
rect 18069 272113 18379 272147
rect 18069 272085 18117 272113
rect 18145 272085 18179 272113
rect 18207 272085 18241 272113
rect 18269 272085 18303 272113
rect 18331 272085 18379 272113
rect 18069 272051 18379 272085
rect 18069 272023 18117 272051
rect 18145 272023 18179 272051
rect 18207 272023 18241 272051
rect 18269 272023 18303 272051
rect 18331 272023 18379 272051
rect 18069 271989 18379 272023
rect 18069 271961 18117 271989
rect 18145 271961 18179 271989
rect 18207 271961 18241 271989
rect 18269 271961 18303 271989
rect 18331 271961 18379 271989
rect 18069 263175 18379 271961
rect 19929 299086 20239 299134
rect 19929 299058 19977 299086
rect 20005 299058 20039 299086
rect 20067 299058 20101 299086
rect 20129 299058 20163 299086
rect 20191 299058 20239 299086
rect 19929 299024 20239 299058
rect 19929 298996 19977 299024
rect 20005 298996 20039 299024
rect 20067 298996 20101 299024
rect 20129 298996 20163 299024
rect 20191 298996 20239 299024
rect 19929 298962 20239 298996
rect 19929 298934 19977 298962
rect 20005 298934 20039 298962
rect 20067 298934 20101 298962
rect 20129 298934 20163 298962
rect 20191 298934 20239 298962
rect 19929 298900 20239 298934
rect 19929 298872 19977 298900
rect 20005 298872 20039 298900
rect 20067 298872 20101 298900
rect 20129 298872 20163 298900
rect 20191 298872 20239 298900
rect 19929 293175 20239 298872
rect 19929 293147 19977 293175
rect 20005 293147 20039 293175
rect 20067 293147 20101 293175
rect 20129 293147 20163 293175
rect 20191 293147 20239 293175
rect 19929 293113 20239 293147
rect 19929 293085 19977 293113
rect 20005 293085 20039 293113
rect 20067 293085 20101 293113
rect 20129 293085 20163 293113
rect 20191 293085 20239 293113
rect 19929 293051 20239 293085
rect 19929 293023 19977 293051
rect 20005 293023 20039 293051
rect 20067 293023 20101 293051
rect 20129 293023 20163 293051
rect 20191 293023 20239 293051
rect 19929 292989 20239 293023
rect 19929 292961 19977 292989
rect 20005 292961 20039 292989
rect 20067 292961 20101 292989
rect 20129 292961 20163 292989
rect 20191 292961 20239 292989
rect 19929 284175 20239 292961
rect 19929 284147 19977 284175
rect 20005 284147 20039 284175
rect 20067 284147 20101 284175
rect 20129 284147 20163 284175
rect 20191 284147 20239 284175
rect 19929 284113 20239 284147
rect 19929 284085 19977 284113
rect 20005 284085 20039 284113
rect 20067 284085 20101 284113
rect 20129 284085 20163 284113
rect 20191 284085 20239 284113
rect 19929 284051 20239 284085
rect 19929 284023 19977 284051
rect 20005 284023 20039 284051
rect 20067 284023 20101 284051
rect 20129 284023 20163 284051
rect 20191 284023 20239 284051
rect 19929 283989 20239 284023
rect 19929 283961 19977 283989
rect 20005 283961 20039 283989
rect 20067 283961 20101 283989
rect 20129 283961 20163 283989
rect 20191 283961 20239 283989
rect 19929 275175 20239 283961
rect 19929 275147 19977 275175
rect 20005 275147 20039 275175
rect 20067 275147 20101 275175
rect 20129 275147 20163 275175
rect 20191 275147 20239 275175
rect 19929 275113 20239 275147
rect 19929 275085 19977 275113
rect 20005 275085 20039 275113
rect 20067 275085 20101 275113
rect 20129 275085 20163 275113
rect 20191 275085 20239 275113
rect 19929 275051 20239 275085
rect 19929 275023 19977 275051
rect 20005 275023 20039 275051
rect 20067 275023 20101 275051
rect 20129 275023 20163 275051
rect 20191 275023 20239 275051
rect 19929 274989 20239 275023
rect 19929 274961 19977 274989
rect 20005 274961 20039 274989
rect 20067 274961 20101 274989
rect 20129 274961 20163 274989
rect 20191 274961 20239 274989
rect 19929 268935 20239 274961
rect 33429 298606 33739 299134
rect 33429 298578 33477 298606
rect 33505 298578 33539 298606
rect 33567 298578 33601 298606
rect 33629 298578 33663 298606
rect 33691 298578 33739 298606
rect 33429 298544 33739 298578
rect 33429 298516 33477 298544
rect 33505 298516 33539 298544
rect 33567 298516 33601 298544
rect 33629 298516 33663 298544
rect 33691 298516 33739 298544
rect 33429 298482 33739 298516
rect 33429 298454 33477 298482
rect 33505 298454 33539 298482
rect 33567 298454 33601 298482
rect 33629 298454 33663 298482
rect 33691 298454 33739 298482
rect 33429 298420 33739 298454
rect 33429 298392 33477 298420
rect 33505 298392 33539 298420
rect 33567 298392 33601 298420
rect 33629 298392 33663 298420
rect 33691 298392 33739 298420
rect 33429 290175 33739 298392
rect 33429 290147 33477 290175
rect 33505 290147 33539 290175
rect 33567 290147 33601 290175
rect 33629 290147 33663 290175
rect 33691 290147 33739 290175
rect 33429 290113 33739 290147
rect 33429 290085 33477 290113
rect 33505 290085 33539 290113
rect 33567 290085 33601 290113
rect 33629 290085 33663 290113
rect 33691 290085 33739 290113
rect 33429 290051 33739 290085
rect 33429 290023 33477 290051
rect 33505 290023 33539 290051
rect 33567 290023 33601 290051
rect 33629 290023 33663 290051
rect 33691 290023 33739 290051
rect 33429 289989 33739 290023
rect 33429 289961 33477 289989
rect 33505 289961 33539 289989
rect 33567 289961 33601 289989
rect 33629 289961 33663 289989
rect 33691 289961 33739 289989
rect 33429 281175 33739 289961
rect 33429 281147 33477 281175
rect 33505 281147 33539 281175
rect 33567 281147 33601 281175
rect 33629 281147 33663 281175
rect 33691 281147 33739 281175
rect 33429 281113 33739 281147
rect 33429 281085 33477 281113
rect 33505 281085 33539 281113
rect 33567 281085 33601 281113
rect 33629 281085 33663 281113
rect 33691 281085 33739 281113
rect 33429 281051 33739 281085
rect 33429 281023 33477 281051
rect 33505 281023 33539 281051
rect 33567 281023 33601 281051
rect 33629 281023 33663 281051
rect 33691 281023 33739 281051
rect 33429 280989 33739 281023
rect 33429 280961 33477 280989
rect 33505 280961 33539 280989
rect 33567 280961 33601 280989
rect 33629 280961 33663 280989
rect 33691 280961 33739 280989
rect 33429 272175 33739 280961
rect 33429 272147 33477 272175
rect 33505 272147 33539 272175
rect 33567 272147 33601 272175
rect 33629 272147 33663 272175
rect 33691 272147 33739 272175
rect 33429 272113 33739 272147
rect 33429 272085 33477 272113
rect 33505 272085 33539 272113
rect 33567 272085 33601 272113
rect 33629 272085 33663 272113
rect 33691 272085 33739 272113
rect 33429 272051 33739 272085
rect 33429 272023 33477 272051
rect 33505 272023 33539 272051
rect 33567 272023 33601 272051
rect 33629 272023 33663 272051
rect 33691 272023 33739 272051
rect 33429 271989 33739 272023
rect 33429 271961 33477 271989
rect 33505 271961 33539 271989
rect 33567 271961 33601 271989
rect 33629 271961 33663 271989
rect 33691 271961 33739 271989
rect 33429 268935 33739 271961
rect 35289 299086 35599 299134
rect 35289 299058 35337 299086
rect 35365 299058 35399 299086
rect 35427 299058 35461 299086
rect 35489 299058 35523 299086
rect 35551 299058 35599 299086
rect 35289 299024 35599 299058
rect 35289 298996 35337 299024
rect 35365 298996 35399 299024
rect 35427 298996 35461 299024
rect 35489 298996 35523 299024
rect 35551 298996 35599 299024
rect 35289 298962 35599 298996
rect 35289 298934 35337 298962
rect 35365 298934 35399 298962
rect 35427 298934 35461 298962
rect 35489 298934 35523 298962
rect 35551 298934 35599 298962
rect 35289 298900 35599 298934
rect 35289 298872 35337 298900
rect 35365 298872 35399 298900
rect 35427 298872 35461 298900
rect 35489 298872 35523 298900
rect 35551 298872 35599 298900
rect 35289 293175 35599 298872
rect 35289 293147 35337 293175
rect 35365 293147 35399 293175
rect 35427 293147 35461 293175
rect 35489 293147 35523 293175
rect 35551 293147 35599 293175
rect 35289 293113 35599 293147
rect 35289 293085 35337 293113
rect 35365 293085 35399 293113
rect 35427 293085 35461 293113
rect 35489 293085 35523 293113
rect 35551 293085 35599 293113
rect 35289 293051 35599 293085
rect 35289 293023 35337 293051
rect 35365 293023 35399 293051
rect 35427 293023 35461 293051
rect 35489 293023 35523 293051
rect 35551 293023 35599 293051
rect 35289 292989 35599 293023
rect 35289 292961 35337 292989
rect 35365 292961 35399 292989
rect 35427 292961 35461 292989
rect 35489 292961 35523 292989
rect 35551 292961 35599 292989
rect 35289 284175 35599 292961
rect 35289 284147 35337 284175
rect 35365 284147 35399 284175
rect 35427 284147 35461 284175
rect 35489 284147 35523 284175
rect 35551 284147 35599 284175
rect 35289 284113 35599 284147
rect 35289 284085 35337 284113
rect 35365 284085 35399 284113
rect 35427 284085 35461 284113
rect 35489 284085 35523 284113
rect 35551 284085 35599 284113
rect 35289 284051 35599 284085
rect 35289 284023 35337 284051
rect 35365 284023 35399 284051
rect 35427 284023 35461 284051
rect 35489 284023 35523 284051
rect 35551 284023 35599 284051
rect 35289 283989 35599 284023
rect 35289 283961 35337 283989
rect 35365 283961 35399 283989
rect 35427 283961 35461 283989
rect 35489 283961 35523 283989
rect 35551 283961 35599 283989
rect 35289 275175 35599 283961
rect 35289 275147 35337 275175
rect 35365 275147 35399 275175
rect 35427 275147 35461 275175
rect 35489 275147 35523 275175
rect 35551 275147 35599 275175
rect 35289 275113 35599 275147
rect 35289 275085 35337 275113
rect 35365 275085 35399 275113
rect 35427 275085 35461 275113
rect 35489 275085 35523 275113
rect 35551 275085 35599 275113
rect 35289 275051 35599 275085
rect 35289 275023 35337 275051
rect 35365 275023 35399 275051
rect 35427 275023 35461 275051
rect 35489 275023 35523 275051
rect 35551 275023 35599 275051
rect 35289 274989 35599 275023
rect 35289 274961 35337 274989
rect 35365 274961 35399 274989
rect 35427 274961 35461 274989
rect 35489 274961 35523 274989
rect 35551 274961 35599 274989
rect 35289 268935 35599 274961
rect 48789 298606 49099 299134
rect 48789 298578 48837 298606
rect 48865 298578 48899 298606
rect 48927 298578 48961 298606
rect 48989 298578 49023 298606
rect 49051 298578 49099 298606
rect 48789 298544 49099 298578
rect 48789 298516 48837 298544
rect 48865 298516 48899 298544
rect 48927 298516 48961 298544
rect 48989 298516 49023 298544
rect 49051 298516 49099 298544
rect 48789 298482 49099 298516
rect 48789 298454 48837 298482
rect 48865 298454 48899 298482
rect 48927 298454 48961 298482
rect 48989 298454 49023 298482
rect 49051 298454 49099 298482
rect 48789 298420 49099 298454
rect 48789 298392 48837 298420
rect 48865 298392 48899 298420
rect 48927 298392 48961 298420
rect 48989 298392 49023 298420
rect 49051 298392 49099 298420
rect 48789 290175 49099 298392
rect 48789 290147 48837 290175
rect 48865 290147 48899 290175
rect 48927 290147 48961 290175
rect 48989 290147 49023 290175
rect 49051 290147 49099 290175
rect 48789 290113 49099 290147
rect 48789 290085 48837 290113
rect 48865 290085 48899 290113
rect 48927 290085 48961 290113
rect 48989 290085 49023 290113
rect 49051 290085 49099 290113
rect 48789 290051 49099 290085
rect 48789 290023 48837 290051
rect 48865 290023 48899 290051
rect 48927 290023 48961 290051
rect 48989 290023 49023 290051
rect 49051 290023 49099 290051
rect 48789 289989 49099 290023
rect 48789 289961 48837 289989
rect 48865 289961 48899 289989
rect 48927 289961 48961 289989
rect 48989 289961 49023 289989
rect 49051 289961 49099 289989
rect 48789 281175 49099 289961
rect 48789 281147 48837 281175
rect 48865 281147 48899 281175
rect 48927 281147 48961 281175
rect 48989 281147 49023 281175
rect 49051 281147 49099 281175
rect 48789 281113 49099 281147
rect 48789 281085 48837 281113
rect 48865 281085 48899 281113
rect 48927 281085 48961 281113
rect 48989 281085 49023 281113
rect 49051 281085 49099 281113
rect 48789 281051 49099 281085
rect 48789 281023 48837 281051
rect 48865 281023 48899 281051
rect 48927 281023 48961 281051
rect 48989 281023 49023 281051
rect 49051 281023 49099 281051
rect 48789 280989 49099 281023
rect 48789 280961 48837 280989
rect 48865 280961 48899 280989
rect 48927 280961 48961 280989
rect 48989 280961 49023 280989
rect 49051 280961 49099 280989
rect 48789 272175 49099 280961
rect 48789 272147 48837 272175
rect 48865 272147 48899 272175
rect 48927 272147 48961 272175
rect 48989 272147 49023 272175
rect 49051 272147 49099 272175
rect 48789 272113 49099 272147
rect 48789 272085 48837 272113
rect 48865 272085 48899 272113
rect 48927 272085 48961 272113
rect 48989 272085 49023 272113
rect 49051 272085 49099 272113
rect 48789 272051 49099 272085
rect 48789 272023 48837 272051
rect 48865 272023 48899 272051
rect 48927 272023 48961 272051
rect 48989 272023 49023 272051
rect 49051 272023 49099 272051
rect 48789 271989 49099 272023
rect 48789 271961 48837 271989
rect 48865 271961 48899 271989
rect 48927 271961 48961 271989
rect 48989 271961 49023 271989
rect 49051 271961 49099 271989
rect 48789 268935 49099 271961
rect 50649 299086 50959 299134
rect 50649 299058 50697 299086
rect 50725 299058 50759 299086
rect 50787 299058 50821 299086
rect 50849 299058 50883 299086
rect 50911 299058 50959 299086
rect 50649 299024 50959 299058
rect 50649 298996 50697 299024
rect 50725 298996 50759 299024
rect 50787 298996 50821 299024
rect 50849 298996 50883 299024
rect 50911 298996 50959 299024
rect 50649 298962 50959 298996
rect 50649 298934 50697 298962
rect 50725 298934 50759 298962
rect 50787 298934 50821 298962
rect 50849 298934 50883 298962
rect 50911 298934 50959 298962
rect 50649 298900 50959 298934
rect 50649 298872 50697 298900
rect 50725 298872 50759 298900
rect 50787 298872 50821 298900
rect 50849 298872 50883 298900
rect 50911 298872 50959 298900
rect 50649 293175 50959 298872
rect 50649 293147 50697 293175
rect 50725 293147 50759 293175
rect 50787 293147 50821 293175
rect 50849 293147 50883 293175
rect 50911 293147 50959 293175
rect 50649 293113 50959 293147
rect 50649 293085 50697 293113
rect 50725 293085 50759 293113
rect 50787 293085 50821 293113
rect 50849 293085 50883 293113
rect 50911 293085 50959 293113
rect 50649 293051 50959 293085
rect 50649 293023 50697 293051
rect 50725 293023 50759 293051
rect 50787 293023 50821 293051
rect 50849 293023 50883 293051
rect 50911 293023 50959 293051
rect 50649 292989 50959 293023
rect 50649 292961 50697 292989
rect 50725 292961 50759 292989
rect 50787 292961 50821 292989
rect 50849 292961 50883 292989
rect 50911 292961 50959 292989
rect 50649 284175 50959 292961
rect 50649 284147 50697 284175
rect 50725 284147 50759 284175
rect 50787 284147 50821 284175
rect 50849 284147 50883 284175
rect 50911 284147 50959 284175
rect 50649 284113 50959 284147
rect 50649 284085 50697 284113
rect 50725 284085 50759 284113
rect 50787 284085 50821 284113
rect 50849 284085 50883 284113
rect 50911 284085 50959 284113
rect 50649 284051 50959 284085
rect 50649 284023 50697 284051
rect 50725 284023 50759 284051
rect 50787 284023 50821 284051
rect 50849 284023 50883 284051
rect 50911 284023 50959 284051
rect 50649 283989 50959 284023
rect 50649 283961 50697 283989
rect 50725 283961 50759 283989
rect 50787 283961 50821 283989
rect 50849 283961 50883 283989
rect 50911 283961 50959 283989
rect 50649 275175 50959 283961
rect 50649 275147 50697 275175
rect 50725 275147 50759 275175
rect 50787 275147 50821 275175
rect 50849 275147 50883 275175
rect 50911 275147 50959 275175
rect 50649 275113 50959 275147
rect 50649 275085 50697 275113
rect 50725 275085 50759 275113
rect 50787 275085 50821 275113
rect 50849 275085 50883 275113
rect 50911 275085 50959 275113
rect 50649 275051 50959 275085
rect 50649 275023 50697 275051
rect 50725 275023 50759 275051
rect 50787 275023 50821 275051
rect 50849 275023 50883 275051
rect 50911 275023 50959 275051
rect 50649 274989 50959 275023
rect 50649 274961 50697 274989
rect 50725 274961 50759 274989
rect 50787 274961 50821 274989
rect 50849 274961 50883 274989
rect 50911 274961 50959 274989
rect 50649 268935 50959 274961
rect 64149 298606 64459 299134
rect 64149 298578 64197 298606
rect 64225 298578 64259 298606
rect 64287 298578 64321 298606
rect 64349 298578 64383 298606
rect 64411 298578 64459 298606
rect 64149 298544 64459 298578
rect 64149 298516 64197 298544
rect 64225 298516 64259 298544
rect 64287 298516 64321 298544
rect 64349 298516 64383 298544
rect 64411 298516 64459 298544
rect 64149 298482 64459 298516
rect 64149 298454 64197 298482
rect 64225 298454 64259 298482
rect 64287 298454 64321 298482
rect 64349 298454 64383 298482
rect 64411 298454 64459 298482
rect 64149 298420 64459 298454
rect 64149 298392 64197 298420
rect 64225 298392 64259 298420
rect 64287 298392 64321 298420
rect 64349 298392 64383 298420
rect 64411 298392 64459 298420
rect 64149 290175 64459 298392
rect 64149 290147 64197 290175
rect 64225 290147 64259 290175
rect 64287 290147 64321 290175
rect 64349 290147 64383 290175
rect 64411 290147 64459 290175
rect 64149 290113 64459 290147
rect 64149 290085 64197 290113
rect 64225 290085 64259 290113
rect 64287 290085 64321 290113
rect 64349 290085 64383 290113
rect 64411 290085 64459 290113
rect 64149 290051 64459 290085
rect 64149 290023 64197 290051
rect 64225 290023 64259 290051
rect 64287 290023 64321 290051
rect 64349 290023 64383 290051
rect 64411 290023 64459 290051
rect 64149 289989 64459 290023
rect 64149 289961 64197 289989
rect 64225 289961 64259 289989
rect 64287 289961 64321 289989
rect 64349 289961 64383 289989
rect 64411 289961 64459 289989
rect 64149 281175 64459 289961
rect 64149 281147 64197 281175
rect 64225 281147 64259 281175
rect 64287 281147 64321 281175
rect 64349 281147 64383 281175
rect 64411 281147 64459 281175
rect 64149 281113 64459 281147
rect 64149 281085 64197 281113
rect 64225 281085 64259 281113
rect 64287 281085 64321 281113
rect 64349 281085 64383 281113
rect 64411 281085 64459 281113
rect 64149 281051 64459 281085
rect 64149 281023 64197 281051
rect 64225 281023 64259 281051
rect 64287 281023 64321 281051
rect 64349 281023 64383 281051
rect 64411 281023 64459 281051
rect 64149 280989 64459 281023
rect 64149 280961 64197 280989
rect 64225 280961 64259 280989
rect 64287 280961 64321 280989
rect 64349 280961 64383 280989
rect 64411 280961 64459 280989
rect 64149 272175 64459 280961
rect 64149 272147 64197 272175
rect 64225 272147 64259 272175
rect 64287 272147 64321 272175
rect 64349 272147 64383 272175
rect 64411 272147 64459 272175
rect 64149 272113 64459 272147
rect 64149 272085 64197 272113
rect 64225 272085 64259 272113
rect 64287 272085 64321 272113
rect 64349 272085 64383 272113
rect 64411 272085 64459 272113
rect 64149 272051 64459 272085
rect 64149 272023 64197 272051
rect 64225 272023 64259 272051
rect 64287 272023 64321 272051
rect 64349 272023 64383 272051
rect 64411 272023 64459 272051
rect 64149 271989 64459 272023
rect 64149 271961 64197 271989
rect 64225 271961 64259 271989
rect 64287 271961 64321 271989
rect 64349 271961 64383 271989
rect 64411 271961 64459 271989
rect 64149 268935 64459 271961
rect 66009 299086 66319 299134
rect 66009 299058 66057 299086
rect 66085 299058 66119 299086
rect 66147 299058 66181 299086
rect 66209 299058 66243 299086
rect 66271 299058 66319 299086
rect 66009 299024 66319 299058
rect 66009 298996 66057 299024
rect 66085 298996 66119 299024
rect 66147 298996 66181 299024
rect 66209 298996 66243 299024
rect 66271 298996 66319 299024
rect 66009 298962 66319 298996
rect 66009 298934 66057 298962
rect 66085 298934 66119 298962
rect 66147 298934 66181 298962
rect 66209 298934 66243 298962
rect 66271 298934 66319 298962
rect 66009 298900 66319 298934
rect 66009 298872 66057 298900
rect 66085 298872 66119 298900
rect 66147 298872 66181 298900
rect 66209 298872 66243 298900
rect 66271 298872 66319 298900
rect 66009 293175 66319 298872
rect 66009 293147 66057 293175
rect 66085 293147 66119 293175
rect 66147 293147 66181 293175
rect 66209 293147 66243 293175
rect 66271 293147 66319 293175
rect 66009 293113 66319 293147
rect 66009 293085 66057 293113
rect 66085 293085 66119 293113
rect 66147 293085 66181 293113
rect 66209 293085 66243 293113
rect 66271 293085 66319 293113
rect 66009 293051 66319 293085
rect 66009 293023 66057 293051
rect 66085 293023 66119 293051
rect 66147 293023 66181 293051
rect 66209 293023 66243 293051
rect 66271 293023 66319 293051
rect 66009 292989 66319 293023
rect 66009 292961 66057 292989
rect 66085 292961 66119 292989
rect 66147 292961 66181 292989
rect 66209 292961 66243 292989
rect 66271 292961 66319 292989
rect 66009 284175 66319 292961
rect 66009 284147 66057 284175
rect 66085 284147 66119 284175
rect 66147 284147 66181 284175
rect 66209 284147 66243 284175
rect 66271 284147 66319 284175
rect 66009 284113 66319 284147
rect 66009 284085 66057 284113
rect 66085 284085 66119 284113
rect 66147 284085 66181 284113
rect 66209 284085 66243 284113
rect 66271 284085 66319 284113
rect 66009 284051 66319 284085
rect 66009 284023 66057 284051
rect 66085 284023 66119 284051
rect 66147 284023 66181 284051
rect 66209 284023 66243 284051
rect 66271 284023 66319 284051
rect 66009 283989 66319 284023
rect 66009 283961 66057 283989
rect 66085 283961 66119 283989
rect 66147 283961 66181 283989
rect 66209 283961 66243 283989
rect 66271 283961 66319 283989
rect 66009 275175 66319 283961
rect 66009 275147 66057 275175
rect 66085 275147 66119 275175
rect 66147 275147 66181 275175
rect 66209 275147 66243 275175
rect 66271 275147 66319 275175
rect 66009 275113 66319 275147
rect 66009 275085 66057 275113
rect 66085 275085 66119 275113
rect 66147 275085 66181 275113
rect 66209 275085 66243 275113
rect 66271 275085 66319 275113
rect 66009 275051 66319 275085
rect 66009 275023 66057 275051
rect 66085 275023 66119 275051
rect 66147 275023 66181 275051
rect 66209 275023 66243 275051
rect 66271 275023 66319 275051
rect 66009 274989 66319 275023
rect 66009 274961 66057 274989
rect 66085 274961 66119 274989
rect 66147 274961 66181 274989
rect 66209 274961 66243 274989
rect 66271 274961 66319 274989
rect 66009 268935 66319 274961
rect 79509 298606 79819 299134
rect 79509 298578 79557 298606
rect 79585 298578 79619 298606
rect 79647 298578 79681 298606
rect 79709 298578 79743 298606
rect 79771 298578 79819 298606
rect 79509 298544 79819 298578
rect 79509 298516 79557 298544
rect 79585 298516 79619 298544
rect 79647 298516 79681 298544
rect 79709 298516 79743 298544
rect 79771 298516 79819 298544
rect 79509 298482 79819 298516
rect 79509 298454 79557 298482
rect 79585 298454 79619 298482
rect 79647 298454 79681 298482
rect 79709 298454 79743 298482
rect 79771 298454 79819 298482
rect 79509 298420 79819 298454
rect 79509 298392 79557 298420
rect 79585 298392 79619 298420
rect 79647 298392 79681 298420
rect 79709 298392 79743 298420
rect 79771 298392 79819 298420
rect 79509 290175 79819 298392
rect 79509 290147 79557 290175
rect 79585 290147 79619 290175
rect 79647 290147 79681 290175
rect 79709 290147 79743 290175
rect 79771 290147 79819 290175
rect 79509 290113 79819 290147
rect 79509 290085 79557 290113
rect 79585 290085 79619 290113
rect 79647 290085 79681 290113
rect 79709 290085 79743 290113
rect 79771 290085 79819 290113
rect 79509 290051 79819 290085
rect 79509 290023 79557 290051
rect 79585 290023 79619 290051
rect 79647 290023 79681 290051
rect 79709 290023 79743 290051
rect 79771 290023 79819 290051
rect 79509 289989 79819 290023
rect 79509 289961 79557 289989
rect 79585 289961 79619 289989
rect 79647 289961 79681 289989
rect 79709 289961 79743 289989
rect 79771 289961 79819 289989
rect 79509 281175 79819 289961
rect 79509 281147 79557 281175
rect 79585 281147 79619 281175
rect 79647 281147 79681 281175
rect 79709 281147 79743 281175
rect 79771 281147 79819 281175
rect 79509 281113 79819 281147
rect 79509 281085 79557 281113
rect 79585 281085 79619 281113
rect 79647 281085 79681 281113
rect 79709 281085 79743 281113
rect 79771 281085 79819 281113
rect 79509 281051 79819 281085
rect 79509 281023 79557 281051
rect 79585 281023 79619 281051
rect 79647 281023 79681 281051
rect 79709 281023 79743 281051
rect 79771 281023 79819 281051
rect 79509 280989 79819 281023
rect 79509 280961 79557 280989
rect 79585 280961 79619 280989
rect 79647 280961 79681 280989
rect 79709 280961 79743 280989
rect 79771 280961 79819 280989
rect 79509 272175 79819 280961
rect 79509 272147 79557 272175
rect 79585 272147 79619 272175
rect 79647 272147 79681 272175
rect 79709 272147 79743 272175
rect 79771 272147 79819 272175
rect 79509 272113 79819 272147
rect 79509 272085 79557 272113
rect 79585 272085 79619 272113
rect 79647 272085 79681 272113
rect 79709 272085 79743 272113
rect 79771 272085 79819 272113
rect 79509 272051 79819 272085
rect 79509 272023 79557 272051
rect 79585 272023 79619 272051
rect 79647 272023 79681 272051
rect 79709 272023 79743 272051
rect 79771 272023 79819 272051
rect 79509 271989 79819 272023
rect 79509 271961 79557 271989
rect 79585 271961 79619 271989
rect 79647 271961 79681 271989
rect 79709 271961 79743 271989
rect 79771 271961 79819 271989
rect 79509 268935 79819 271961
rect 81369 299086 81679 299134
rect 81369 299058 81417 299086
rect 81445 299058 81479 299086
rect 81507 299058 81541 299086
rect 81569 299058 81603 299086
rect 81631 299058 81679 299086
rect 81369 299024 81679 299058
rect 81369 298996 81417 299024
rect 81445 298996 81479 299024
rect 81507 298996 81541 299024
rect 81569 298996 81603 299024
rect 81631 298996 81679 299024
rect 81369 298962 81679 298996
rect 81369 298934 81417 298962
rect 81445 298934 81479 298962
rect 81507 298934 81541 298962
rect 81569 298934 81603 298962
rect 81631 298934 81679 298962
rect 81369 298900 81679 298934
rect 81369 298872 81417 298900
rect 81445 298872 81479 298900
rect 81507 298872 81541 298900
rect 81569 298872 81603 298900
rect 81631 298872 81679 298900
rect 81369 293175 81679 298872
rect 81369 293147 81417 293175
rect 81445 293147 81479 293175
rect 81507 293147 81541 293175
rect 81569 293147 81603 293175
rect 81631 293147 81679 293175
rect 81369 293113 81679 293147
rect 81369 293085 81417 293113
rect 81445 293085 81479 293113
rect 81507 293085 81541 293113
rect 81569 293085 81603 293113
rect 81631 293085 81679 293113
rect 81369 293051 81679 293085
rect 81369 293023 81417 293051
rect 81445 293023 81479 293051
rect 81507 293023 81541 293051
rect 81569 293023 81603 293051
rect 81631 293023 81679 293051
rect 81369 292989 81679 293023
rect 81369 292961 81417 292989
rect 81445 292961 81479 292989
rect 81507 292961 81541 292989
rect 81569 292961 81603 292989
rect 81631 292961 81679 292989
rect 81369 284175 81679 292961
rect 81369 284147 81417 284175
rect 81445 284147 81479 284175
rect 81507 284147 81541 284175
rect 81569 284147 81603 284175
rect 81631 284147 81679 284175
rect 81369 284113 81679 284147
rect 81369 284085 81417 284113
rect 81445 284085 81479 284113
rect 81507 284085 81541 284113
rect 81569 284085 81603 284113
rect 81631 284085 81679 284113
rect 81369 284051 81679 284085
rect 81369 284023 81417 284051
rect 81445 284023 81479 284051
rect 81507 284023 81541 284051
rect 81569 284023 81603 284051
rect 81631 284023 81679 284051
rect 81369 283989 81679 284023
rect 81369 283961 81417 283989
rect 81445 283961 81479 283989
rect 81507 283961 81541 283989
rect 81569 283961 81603 283989
rect 81631 283961 81679 283989
rect 81369 275175 81679 283961
rect 81369 275147 81417 275175
rect 81445 275147 81479 275175
rect 81507 275147 81541 275175
rect 81569 275147 81603 275175
rect 81631 275147 81679 275175
rect 81369 275113 81679 275147
rect 81369 275085 81417 275113
rect 81445 275085 81479 275113
rect 81507 275085 81541 275113
rect 81569 275085 81603 275113
rect 81631 275085 81679 275113
rect 81369 275051 81679 275085
rect 81369 275023 81417 275051
rect 81445 275023 81479 275051
rect 81507 275023 81541 275051
rect 81569 275023 81603 275051
rect 81631 275023 81679 275051
rect 81369 274989 81679 275023
rect 81369 274961 81417 274989
rect 81445 274961 81479 274989
rect 81507 274961 81541 274989
rect 81569 274961 81603 274989
rect 81631 274961 81679 274989
rect 81369 268935 81679 274961
rect 94869 298606 95179 299134
rect 94869 298578 94917 298606
rect 94945 298578 94979 298606
rect 95007 298578 95041 298606
rect 95069 298578 95103 298606
rect 95131 298578 95179 298606
rect 94869 298544 95179 298578
rect 94869 298516 94917 298544
rect 94945 298516 94979 298544
rect 95007 298516 95041 298544
rect 95069 298516 95103 298544
rect 95131 298516 95179 298544
rect 94869 298482 95179 298516
rect 94869 298454 94917 298482
rect 94945 298454 94979 298482
rect 95007 298454 95041 298482
rect 95069 298454 95103 298482
rect 95131 298454 95179 298482
rect 94869 298420 95179 298454
rect 94869 298392 94917 298420
rect 94945 298392 94979 298420
rect 95007 298392 95041 298420
rect 95069 298392 95103 298420
rect 95131 298392 95179 298420
rect 94869 290175 95179 298392
rect 94869 290147 94917 290175
rect 94945 290147 94979 290175
rect 95007 290147 95041 290175
rect 95069 290147 95103 290175
rect 95131 290147 95179 290175
rect 94869 290113 95179 290147
rect 94869 290085 94917 290113
rect 94945 290085 94979 290113
rect 95007 290085 95041 290113
rect 95069 290085 95103 290113
rect 95131 290085 95179 290113
rect 94869 290051 95179 290085
rect 94869 290023 94917 290051
rect 94945 290023 94979 290051
rect 95007 290023 95041 290051
rect 95069 290023 95103 290051
rect 95131 290023 95179 290051
rect 94869 289989 95179 290023
rect 94869 289961 94917 289989
rect 94945 289961 94979 289989
rect 95007 289961 95041 289989
rect 95069 289961 95103 289989
rect 95131 289961 95179 289989
rect 94869 281175 95179 289961
rect 94869 281147 94917 281175
rect 94945 281147 94979 281175
rect 95007 281147 95041 281175
rect 95069 281147 95103 281175
rect 95131 281147 95179 281175
rect 94869 281113 95179 281147
rect 94869 281085 94917 281113
rect 94945 281085 94979 281113
rect 95007 281085 95041 281113
rect 95069 281085 95103 281113
rect 95131 281085 95179 281113
rect 94869 281051 95179 281085
rect 94869 281023 94917 281051
rect 94945 281023 94979 281051
rect 95007 281023 95041 281051
rect 95069 281023 95103 281051
rect 95131 281023 95179 281051
rect 94869 280989 95179 281023
rect 94869 280961 94917 280989
rect 94945 280961 94979 280989
rect 95007 280961 95041 280989
rect 95069 280961 95103 280989
rect 95131 280961 95179 280989
rect 94869 272175 95179 280961
rect 94869 272147 94917 272175
rect 94945 272147 94979 272175
rect 95007 272147 95041 272175
rect 95069 272147 95103 272175
rect 95131 272147 95179 272175
rect 94869 272113 95179 272147
rect 94869 272085 94917 272113
rect 94945 272085 94979 272113
rect 95007 272085 95041 272113
rect 95069 272085 95103 272113
rect 95131 272085 95179 272113
rect 94869 272051 95179 272085
rect 94869 272023 94917 272051
rect 94945 272023 94979 272051
rect 95007 272023 95041 272051
rect 95069 272023 95103 272051
rect 95131 272023 95179 272051
rect 94869 271989 95179 272023
rect 94869 271961 94917 271989
rect 94945 271961 94979 271989
rect 95007 271961 95041 271989
rect 95069 271961 95103 271989
rect 95131 271961 95179 271989
rect 29904 266175 30064 266192
rect 29904 266147 29939 266175
rect 29967 266147 30001 266175
rect 30029 266147 30064 266175
rect 29904 266113 30064 266147
rect 29904 266085 29939 266113
rect 29967 266085 30001 266113
rect 30029 266085 30064 266113
rect 29904 266051 30064 266085
rect 29904 266023 29939 266051
rect 29967 266023 30001 266051
rect 30029 266023 30064 266051
rect 29904 265989 30064 266023
rect 29904 265961 29939 265989
rect 29967 265961 30001 265989
rect 30029 265961 30064 265989
rect 29904 265944 30064 265961
rect 45264 266175 45424 266192
rect 45264 266147 45299 266175
rect 45327 266147 45361 266175
rect 45389 266147 45424 266175
rect 45264 266113 45424 266147
rect 45264 266085 45299 266113
rect 45327 266085 45361 266113
rect 45389 266085 45424 266113
rect 45264 266051 45424 266085
rect 45264 266023 45299 266051
rect 45327 266023 45361 266051
rect 45389 266023 45424 266051
rect 45264 265989 45424 266023
rect 45264 265961 45299 265989
rect 45327 265961 45361 265989
rect 45389 265961 45424 265989
rect 45264 265944 45424 265961
rect 60624 266175 60784 266192
rect 60624 266147 60659 266175
rect 60687 266147 60721 266175
rect 60749 266147 60784 266175
rect 60624 266113 60784 266147
rect 60624 266085 60659 266113
rect 60687 266085 60721 266113
rect 60749 266085 60784 266113
rect 60624 266051 60784 266085
rect 60624 266023 60659 266051
rect 60687 266023 60721 266051
rect 60749 266023 60784 266051
rect 60624 265989 60784 266023
rect 60624 265961 60659 265989
rect 60687 265961 60721 265989
rect 60749 265961 60784 265989
rect 60624 265944 60784 265961
rect 75984 266175 76144 266192
rect 75984 266147 76019 266175
rect 76047 266147 76081 266175
rect 76109 266147 76144 266175
rect 75984 266113 76144 266147
rect 75984 266085 76019 266113
rect 76047 266085 76081 266113
rect 76109 266085 76144 266113
rect 75984 266051 76144 266085
rect 75984 266023 76019 266051
rect 76047 266023 76081 266051
rect 76109 266023 76144 266051
rect 75984 265989 76144 266023
rect 75984 265961 76019 265989
rect 76047 265961 76081 265989
rect 76109 265961 76144 265989
rect 75984 265944 76144 265961
rect 18069 263147 18117 263175
rect 18145 263147 18179 263175
rect 18207 263147 18241 263175
rect 18269 263147 18303 263175
rect 18331 263147 18379 263175
rect 18069 263113 18379 263147
rect 18069 263085 18117 263113
rect 18145 263085 18179 263113
rect 18207 263085 18241 263113
rect 18269 263085 18303 263113
rect 18331 263085 18379 263113
rect 18069 263051 18379 263085
rect 18069 263023 18117 263051
rect 18145 263023 18179 263051
rect 18207 263023 18241 263051
rect 18269 263023 18303 263051
rect 18331 263023 18379 263051
rect 18069 262989 18379 263023
rect 18069 262961 18117 262989
rect 18145 262961 18179 262989
rect 18207 262961 18241 262989
rect 18269 262961 18303 262989
rect 18331 262961 18379 262989
rect 5446 154961 5474 154966
rect 5502 258314 5530 258319
rect 5502 153314 5530 258286
rect 18069 254175 18379 262961
rect 22224 263175 22384 263192
rect 22224 263147 22259 263175
rect 22287 263147 22321 263175
rect 22349 263147 22384 263175
rect 22224 263113 22384 263147
rect 22224 263085 22259 263113
rect 22287 263085 22321 263113
rect 22349 263085 22384 263113
rect 22224 263051 22384 263085
rect 22224 263023 22259 263051
rect 22287 263023 22321 263051
rect 22349 263023 22384 263051
rect 22224 262989 22384 263023
rect 22224 262961 22259 262989
rect 22287 262961 22321 262989
rect 22349 262961 22384 262989
rect 22224 262944 22384 262961
rect 37584 263175 37744 263192
rect 37584 263147 37619 263175
rect 37647 263147 37681 263175
rect 37709 263147 37744 263175
rect 37584 263113 37744 263147
rect 37584 263085 37619 263113
rect 37647 263085 37681 263113
rect 37709 263085 37744 263113
rect 37584 263051 37744 263085
rect 37584 263023 37619 263051
rect 37647 263023 37681 263051
rect 37709 263023 37744 263051
rect 37584 262989 37744 263023
rect 37584 262961 37619 262989
rect 37647 262961 37681 262989
rect 37709 262961 37744 262989
rect 37584 262944 37744 262961
rect 52944 263175 53104 263192
rect 52944 263147 52979 263175
rect 53007 263147 53041 263175
rect 53069 263147 53104 263175
rect 52944 263113 53104 263147
rect 52944 263085 52979 263113
rect 53007 263085 53041 263113
rect 53069 263085 53104 263113
rect 52944 263051 53104 263085
rect 52944 263023 52979 263051
rect 53007 263023 53041 263051
rect 53069 263023 53104 263051
rect 52944 262989 53104 263023
rect 52944 262961 52979 262989
rect 53007 262961 53041 262989
rect 53069 262961 53104 262989
rect 52944 262944 53104 262961
rect 68304 263175 68464 263192
rect 68304 263147 68339 263175
rect 68367 263147 68401 263175
rect 68429 263147 68464 263175
rect 68304 263113 68464 263147
rect 68304 263085 68339 263113
rect 68367 263085 68401 263113
rect 68429 263085 68464 263113
rect 68304 263051 68464 263085
rect 68304 263023 68339 263051
rect 68367 263023 68401 263051
rect 68429 263023 68464 263051
rect 68304 262989 68464 263023
rect 68304 262961 68339 262989
rect 68367 262961 68401 262989
rect 68429 262961 68464 262989
rect 68304 262944 68464 262961
rect 83664 263175 83824 263192
rect 83664 263147 83699 263175
rect 83727 263147 83761 263175
rect 83789 263147 83824 263175
rect 83664 263113 83824 263147
rect 83664 263085 83699 263113
rect 83727 263085 83761 263113
rect 83789 263085 83824 263113
rect 83664 263051 83824 263085
rect 83664 263023 83699 263051
rect 83727 263023 83761 263051
rect 83789 263023 83824 263051
rect 83664 262989 83824 263023
rect 83664 262961 83699 262989
rect 83727 262961 83761 262989
rect 83789 262961 83824 262989
rect 83664 262944 83824 262961
rect 94869 263175 95179 271961
rect 94869 263147 94917 263175
rect 94945 263147 94979 263175
rect 95007 263147 95041 263175
rect 95069 263147 95103 263175
rect 95131 263147 95179 263175
rect 94869 263113 95179 263147
rect 94869 263085 94917 263113
rect 94945 263085 94979 263113
rect 95007 263085 95041 263113
rect 95069 263085 95103 263113
rect 95131 263085 95179 263113
rect 94869 263051 95179 263085
rect 94869 263023 94917 263051
rect 94945 263023 94979 263051
rect 95007 263023 95041 263051
rect 95069 263023 95103 263051
rect 95131 263023 95179 263051
rect 94869 262989 95179 263023
rect 94869 262961 94917 262989
rect 94945 262961 94979 262989
rect 95007 262961 95041 262989
rect 95069 262961 95103 262989
rect 95131 262961 95179 262989
rect 29904 257175 30064 257192
rect 29904 257147 29939 257175
rect 29967 257147 30001 257175
rect 30029 257147 30064 257175
rect 29904 257113 30064 257147
rect 29904 257085 29939 257113
rect 29967 257085 30001 257113
rect 30029 257085 30064 257113
rect 29904 257051 30064 257085
rect 29904 257023 29939 257051
rect 29967 257023 30001 257051
rect 30029 257023 30064 257051
rect 29904 256989 30064 257023
rect 29904 256961 29939 256989
rect 29967 256961 30001 256989
rect 30029 256961 30064 256989
rect 29904 256944 30064 256961
rect 45264 257175 45424 257192
rect 45264 257147 45299 257175
rect 45327 257147 45361 257175
rect 45389 257147 45424 257175
rect 45264 257113 45424 257147
rect 45264 257085 45299 257113
rect 45327 257085 45361 257113
rect 45389 257085 45424 257113
rect 45264 257051 45424 257085
rect 45264 257023 45299 257051
rect 45327 257023 45361 257051
rect 45389 257023 45424 257051
rect 45264 256989 45424 257023
rect 45264 256961 45299 256989
rect 45327 256961 45361 256989
rect 45389 256961 45424 256989
rect 45264 256944 45424 256961
rect 60624 257175 60784 257192
rect 60624 257147 60659 257175
rect 60687 257147 60721 257175
rect 60749 257147 60784 257175
rect 60624 257113 60784 257147
rect 60624 257085 60659 257113
rect 60687 257085 60721 257113
rect 60749 257085 60784 257113
rect 60624 257051 60784 257085
rect 60624 257023 60659 257051
rect 60687 257023 60721 257051
rect 60749 257023 60784 257051
rect 60624 256989 60784 257023
rect 60624 256961 60659 256989
rect 60687 256961 60721 256989
rect 60749 256961 60784 256989
rect 60624 256944 60784 256961
rect 75984 257175 76144 257192
rect 75984 257147 76019 257175
rect 76047 257147 76081 257175
rect 76109 257147 76144 257175
rect 75984 257113 76144 257147
rect 75984 257085 76019 257113
rect 76047 257085 76081 257113
rect 76109 257085 76144 257113
rect 75984 257051 76144 257085
rect 75984 257023 76019 257051
rect 76047 257023 76081 257051
rect 76109 257023 76144 257051
rect 75984 256989 76144 257023
rect 75984 256961 76019 256989
rect 76047 256961 76081 256989
rect 76109 256961 76144 256989
rect 75984 256944 76144 256961
rect 18069 254147 18117 254175
rect 18145 254147 18179 254175
rect 18207 254147 18241 254175
rect 18269 254147 18303 254175
rect 18331 254147 18379 254175
rect 18069 254113 18379 254147
rect 18069 254085 18117 254113
rect 18145 254085 18179 254113
rect 18207 254085 18241 254113
rect 18269 254085 18303 254113
rect 18331 254085 18379 254113
rect 18069 254051 18379 254085
rect 18069 254023 18117 254051
rect 18145 254023 18179 254051
rect 18207 254023 18241 254051
rect 18269 254023 18303 254051
rect 18331 254023 18379 254051
rect 18069 253989 18379 254023
rect 18069 253961 18117 253989
rect 18145 253961 18179 253989
rect 18207 253961 18241 253989
rect 18269 253961 18303 253989
rect 18331 253961 18379 253989
rect 18069 245175 18379 253961
rect 22224 254175 22384 254192
rect 22224 254147 22259 254175
rect 22287 254147 22321 254175
rect 22349 254147 22384 254175
rect 22224 254113 22384 254147
rect 22224 254085 22259 254113
rect 22287 254085 22321 254113
rect 22349 254085 22384 254113
rect 22224 254051 22384 254085
rect 22224 254023 22259 254051
rect 22287 254023 22321 254051
rect 22349 254023 22384 254051
rect 22224 253989 22384 254023
rect 22224 253961 22259 253989
rect 22287 253961 22321 253989
rect 22349 253961 22384 253989
rect 22224 253944 22384 253961
rect 37584 254175 37744 254192
rect 37584 254147 37619 254175
rect 37647 254147 37681 254175
rect 37709 254147 37744 254175
rect 37584 254113 37744 254147
rect 37584 254085 37619 254113
rect 37647 254085 37681 254113
rect 37709 254085 37744 254113
rect 37584 254051 37744 254085
rect 37584 254023 37619 254051
rect 37647 254023 37681 254051
rect 37709 254023 37744 254051
rect 37584 253989 37744 254023
rect 37584 253961 37619 253989
rect 37647 253961 37681 253989
rect 37709 253961 37744 253989
rect 37584 253944 37744 253961
rect 52944 254175 53104 254192
rect 52944 254147 52979 254175
rect 53007 254147 53041 254175
rect 53069 254147 53104 254175
rect 52944 254113 53104 254147
rect 52944 254085 52979 254113
rect 53007 254085 53041 254113
rect 53069 254085 53104 254113
rect 52944 254051 53104 254085
rect 52944 254023 52979 254051
rect 53007 254023 53041 254051
rect 53069 254023 53104 254051
rect 52944 253989 53104 254023
rect 52944 253961 52979 253989
rect 53007 253961 53041 253989
rect 53069 253961 53104 253989
rect 52944 253944 53104 253961
rect 68304 254175 68464 254192
rect 68304 254147 68339 254175
rect 68367 254147 68401 254175
rect 68429 254147 68464 254175
rect 68304 254113 68464 254147
rect 68304 254085 68339 254113
rect 68367 254085 68401 254113
rect 68429 254085 68464 254113
rect 68304 254051 68464 254085
rect 68304 254023 68339 254051
rect 68367 254023 68401 254051
rect 68429 254023 68464 254051
rect 68304 253989 68464 254023
rect 68304 253961 68339 253989
rect 68367 253961 68401 253989
rect 68429 253961 68464 253989
rect 68304 253944 68464 253961
rect 83664 254175 83824 254192
rect 83664 254147 83699 254175
rect 83727 254147 83761 254175
rect 83789 254147 83824 254175
rect 83664 254113 83824 254147
rect 83664 254085 83699 254113
rect 83727 254085 83761 254113
rect 83789 254085 83824 254113
rect 83664 254051 83824 254085
rect 83664 254023 83699 254051
rect 83727 254023 83761 254051
rect 83789 254023 83824 254051
rect 83664 253989 83824 254023
rect 83664 253961 83699 253989
rect 83727 253961 83761 253989
rect 83789 253961 83824 253989
rect 83664 253944 83824 253961
rect 94869 254175 95179 262961
rect 94869 254147 94917 254175
rect 94945 254147 94979 254175
rect 95007 254147 95041 254175
rect 95069 254147 95103 254175
rect 95131 254147 95179 254175
rect 94869 254113 95179 254147
rect 94869 254085 94917 254113
rect 94945 254085 94979 254113
rect 95007 254085 95041 254113
rect 95069 254085 95103 254113
rect 95131 254085 95179 254113
rect 94869 254051 95179 254085
rect 94869 254023 94917 254051
rect 94945 254023 94979 254051
rect 95007 254023 95041 254051
rect 95069 254023 95103 254051
rect 95131 254023 95179 254051
rect 94869 253989 95179 254023
rect 94869 253961 94917 253989
rect 94945 253961 94979 253989
rect 95007 253961 95041 253989
rect 95069 253961 95103 253989
rect 95131 253961 95179 253989
rect 29904 248175 30064 248192
rect 29904 248147 29939 248175
rect 29967 248147 30001 248175
rect 30029 248147 30064 248175
rect 29904 248113 30064 248147
rect 29904 248085 29939 248113
rect 29967 248085 30001 248113
rect 30029 248085 30064 248113
rect 29904 248051 30064 248085
rect 29904 248023 29939 248051
rect 29967 248023 30001 248051
rect 30029 248023 30064 248051
rect 29904 247989 30064 248023
rect 29904 247961 29939 247989
rect 29967 247961 30001 247989
rect 30029 247961 30064 247989
rect 29904 247944 30064 247961
rect 45264 248175 45424 248192
rect 45264 248147 45299 248175
rect 45327 248147 45361 248175
rect 45389 248147 45424 248175
rect 45264 248113 45424 248147
rect 45264 248085 45299 248113
rect 45327 248085 45361 248113
rect 45389 248085 45424 248113
rect 45264 248051 45424 248085
rect 45264 248023 45299 248051
rect 45327 248023 45361 248051
rect 45389 248023 45424 248051
rect 45264 247989 45424 248023
rect 45264 247961 45299 247989
rect 45327 247961 45361 247989
rect 45389 247961 45424 247989
rect 45264 247944 45424 247961
rect 60624 248175 60784 248192
rect 60624 248147 60659 248175
rect 60687 248147 60721 248175
rect 60749 248147 60784 248175
rect 60624 248113 60784 248147
rect 60624 248085 60659 248113
rect 60687 248085 60721 248113
rect 60749 248085 60784 248113
rect 60624 248051 60784 248085
rect 60624 248023 60659 248051
rect 60687 248023 60721 248051
rect 60749 248023 60784 248051
rect 60624 247989 60784 248023
rect 60624 247961 60659 247989
rect 60687 247961 60721 247989
rect 60749 247961 60784 247989
rect 60624 247944 60784 247961
rect 75984 248175 76144 248192
rect 75984 248147 76019 248175
rect 76047 248147 76081 248175
rect 76109 248147 76144 248175
rect 75984 248113 76144 248147
rect 75984 248085 76019 248113
rect 76047 248085 76081 248113
rect 76109 248085 76144 248113
rect 75984 248051 76144 248085
rect 75984 248023 76019 248051
rect 76047 248023 76081 248051
rect 76109 248023 76144 248051
rect 75984 247989 76144 248023
rect 75984 247961 76019 247989
rect 76047 247961 76081 247989
rect 76109 247961 76144 247989
rect 75984 247944 76144 247961
rect 18069 245147 18117 245175
rect 18145 245147 18179 245175
rect 18207 245147 18241 245175
rect 18269 245147 18303 245175
rect 18331 245147 18379 245175
rect 18069 245113 18379 245147
rect 18069 245085 18117 245113
rect 18145 245085 18179 245113
rect 18207 245085 18241 245113
rect 18269 245085 18303 245113
rect 18331 245085 18379 245113
rect 18069 245051 18379 245085
rect 18069 245023 18117 245051
rect 18145 245023 18179 245051
rect 18207 245023 18241 245051
rect 18269 245023 18303 245051
rect 18331 245023 18379 245051
rect 18069 244989 18379 245023
rect 18069 244961 18117 244989
rect 18145 244961 18179 244989
rect 18207 244961 18241 244989
rect 18269 244961 18303 244989
rect 18331 244961 18379 244989
rect 5502 153281 5530 153286
rect 5558 237146 5586 237151
rect 5558 151634 5586 237118
rect 18069 236175 18379 244961
rect 22224 245175 22384 245192
rect 22224 245147 22259 245175
rect 22287 245147 22321 245175
rect 22349 245147 22384 245175
rect 22224 245113 22384 245147
rect 22224 245085 22259 245113
rect 22287 245085 22321 245113
rect 22349 245085 22384 245113
rect 22224 245051 22384 245085
rect 22224 245023 22259 245051
rect 22287 245023 22321 245051
rect 22349 245023 22384 245051
rect 22224 244989 22384 245023
rect 22224 244961 22259 244989
rect 22287 244961 22321 244989
rect 22349 244961 22384 244989
rect 22224 244944 22384 244961
rect 37584 245175 37744 245192
rect 37584 245147 37619 245175
rect 37647 245147 37681 245175
rect 37709 245147 37744 245175
rect 37584 245113 37744 245147
rect 37584 245085 37619 245113
rect 37647 245085 37681 245113
rect 37709 245085 37744 245113
rect 37584 245051 37744 245085
rect 37584 245023 37619 245051
rect 37647 245023 37681 245051
rect 37709 245023 37744 245051
rect 37584 244989 37744 245023
rect 37584 244961 37619 244989
rect 37647 244961 37681 244989
rect 37709 244961 37744 244989
rect 37584 244944 37744 244961
rect 52944 245175 53104 245192
rect 52944 245147 52979 245175
rect 53007 245147 53041 245175
rect 53069 245147 53104 245175
rect 52944 245113 53104 245147
rect 52944 245085 52979 245113
rect 53007 245085 53041 245113
rect 53069 245085 53104 245113
rect 52944 245051 53104 245085
rect 52944 245023 52979 245051
rect 53007 245023 53041 245051
rect 53069 245023 53104 245051
rect 52944 244989 53104 245023
rect 52944 244961 52979 244989
rect 53007 244961 53041 244989
rect 53069 244961 53104 244989
rect 52944 244944 53104 244961
rect 68304 245175 68464 245192
rect 68304 245147 68339 245175
rect 68367 245147 68401 245175
rect 68429 245147 68464 245175
rect 68304 245113 68464 245147
rect 68304 245085 68339 245113
rect 68367 245085 68401 245113
rect 68429 245085 68464 245113
rect 68304 245051 68464 245085
rect 68304 245023 68339 245051
rect 68367 245023 68401 245051
rect 68429 245023 68464 245051
rect 68304 244989 68464 245023
rect 68304 244961 68339 244989
rect 68367 244961 68401 244989
rect 68429 244961 68464 244989
rect 68304 244944 68464 244961
rect 83664 245175 83824 245192
rect 83664 245147 83699 245175
rect 83727 245147 83761 245175
rect 83789 245147 83824 245175
rect 83664 245113 83824 245147
rect 83664 245085 83699 245113
rect 83727 245085 83761 245113
rect 83789 245085 83824 245113
rect 83664 245051 83824 245085
rect 83664 245023 83699 245051
rect 83727 245023 83761 245051
rect 83789 245023 83824 245051
rect 83664 244989 83824 245023
rect 83664 244961 83699 244989
rect 83727 244961 83761 244989
rect 83789 244961 83824 244989
rect 83664 244944 83824 244961
rect 94869 245175 95179 253961
rect 94869 245147 94917 245175
rect 94945 245147 94979 245175
rect 95007 245147 95041 245175
rect 95069 245147 95103 245175
rect 95131 245147 95179 245175
rect 94869 245113 95179 245147
rect 94869 245085 94917 245113
rect 94945 245085 94979 245113
rect 95007 245085 95041 245113
rect 95069 245085 95103 245113
rect 95131 245085 95179 245113
rect 94869 245051 95179 245085
rect 94869 245023 94917 245051
rect 94945 245023 94979 245051
rect 95007 245023 95041 245051
rect 95069 245023 95103 245051
rect 95131 245023 95179 245051
rect 94869 244989 95179 245023
rect 94869 244961 94917 244989
rect 94945 244961 94979 244989
rect 95007 244961 95041 244989
rect 95069 244961 95103 244989
rect 95131 244961 95179 244989
rect 29904 239175 30064 239192
rect 29904 239147 29939 239175
rect 29967 239147 30001 239175
rect 30029 239147 30064 239175
rect 29904 239113 30064 239147
rect 29904 239085 29939 239113
rect 29967 239085 30001 239113
rect 30029 239085 30064 239113
rect 29904 239051 30064 239085
rect 29904 239023 29939 239051
rect 29967 239023 30001 239051
rect 30029 239023 30064 239051
rect 29904 238989 30064 239023
rect 29904 238961 29939 238989
rect 29967 238961 30001 238989
rect 30029 238961 30064 238989
rect 29904 238944 30064 238961
rect 45264 239175 45424 239192
rect 45264 239147 45299 239175
rect 45327 239147 45361 239175
rect 45389 239147 45424 239175
rect 45264 239113 45424 239147
rect 45264 239085 45299 239113
rect 45327 239085 45361 239113
rect 45389 239085 45424 239113
rect 45264 239051 45424 239085
rect 45264 239023 45299 239051
rect 45327 239023 45361 239051
rect 45389 239023 45424 239051
rect 45264 238989 45424 239023
rect 45264 238961 45299 238989
rect 45327 238961 45361 238989
rect 45389 238961 45424 238989
rect 45264 238944 45424 238961
rect 60624 239175 60784 239192
rect 60624 239147 60659 239175
rect 60687 239147 60721 239175
rect 60749 239147 60784 239175
rect 60624 239113 60784 239147
rect 60624 239085 60659 239113
rect 60687 239085 60721 239113
rect 60749 239085 60784 239113
rect 60624 239051 60784 239085
rect 60624 239023 60659 239051
rect 60687 239023 60721 239051
rect 60749 239023 60784 239051
rect 60624 238989 60784 239023
rect 60624 238961 60659 238989
rect 60687 238961 60721 238989
rect 60749 238961 60784 238989
rect 60624 238944 60784 238961
rect 75984 239175 76144 239192
rect 75984 239147 76019 239175
rect 76047 239147 76081 239175
rect 76109 239147 76144 239175
rect 75984 239113 76144 239147
rect 75984 239085 76019 239113
rect 76047 239085 76081 239113
rect 76109 239085 76144 239113
rect 75984 239051 76144 239085
rect 75984 239023 76019 239051
rect 76047 239023 76081 239051
rect 76109 239023 76144 239051
rect 75984 238989 76144 239023
rect 75984 238961 76019 238989
rect 76047 238961 76081 238989
rect 76109 238961 76144 238989
rect 75984 238944 76144 238961
rect 18069 236147 18117 236175
rect 18145 236147 18179 236175
rect 18207 236147 18241 236175
rect 18269 236147 18303 236175
rect 18331 236147 18379 236175
rect 18069 236113 18379 236147
rect 18069 236085 18117 236113
rect 18145 236085 18179 236113
rect 18207 236085 18241 236113
rect 18269 236085 18303 236113
rect 18331 236085 18379 236113
rect 18069 236051 18379 236085
rect 18069 236023 18117 236051
rect 18145 236023 18179 236051
rect 18207 236023 18241 236051
rect 18269 236023 18303 236051
rect 18331 236023 18379 236051
rect 18069 235989 18379 236023
rect 18069 235961 18117 235989
rect 18145 235961 18179 235989
rect 18207 235961 18241 235989
rect 18269 235961 18303 235989
rect 18331 235961 18379 235989
rect 18069 227175 18379 235961
rect 22224 236175 22384 236192
rect 22224 236147 22259 236175
rect 22287 236147 22321 236175
rect 22349 236147 22384 236175
rect 22224 236113 22384 236147
rect 22224 236085 22259 236113
rect 22287 236085 22321 236113
rect 22349 236085 22384 236113
rect 22224 236051 22384 236085
rect 22224 236023 22259 236051
rect 22287 236023 22321 236051
rect 22349 236023 22384 236051
rect 22224 235989 22384 236023
rect 22224 235961 22259 235989
rect 22287 235961 22321 235989
rect 22349 235961 22384 235989
rect 22224 235944 22384 235961
rect 37584 236175 37744 236192
rect 37584 236147 37619 236175
rect 37647 236147 37681 236175
rect 37709 236147 37744 236175
rect 37584 236113 37744 236147
rect 37584 236085 37619 236113
rect 37647 236085 37681 236113
rect 37709 236085 37744 236113
rect 37584 236051 37744 236085
rect 37584 236023 37619 236051
rect 37647 236023 37681 236051
rect 37709 236023 37744 236051
rect 37584 235989 37744 236023
rect 37584 235961 37619 235989
rect 37647 235961 37681 235989
rect 37709 235961 37744 235989
rect 37584 235944 37744 235961
rect 52944 236175 53104 236192
rect 52944 236147 52979 236175
rect 53007 236147 53041 236175
rect 53069 236147 53104 236175
rect 52944 236113 53104 236147
rect 52944 236085 52979 236113
rect 53007 236085 53041 236113
rect 53069 236085 53104 236113
rect 52944 236051 53104 236085
rect 52944 236023 52979 236051
rect 53007 236023 53041 236051
rect 53069 236023 53104 236051
rect 52944 235989 53104 236023
rect 52944 235961 52979 235989
rect 53007 235961 53041 235989
rect 53069 235961 53104 235989
rect 52944 235944 53104 235961
rect 68304 236175 68464 236192
rect 68304 236147 68339 236175
rect 68367 236147 68401 236175
rect 68429 236147 68464 236175
rect 68304 236113 68464 236147
rect 68304 236085 68339 236113
rect 68367 236085 68401 236113
rect 68429 236085 68464 236113
rect 68304 236051 68464 236085
rect 68304 236023 68339 236051
rect 68367 236023 68401 236051
rect 68429 236023 68464 236051
rect 68304 235989 68464 236023
rect 68304 235961 68339 235989
rect 68367 235961 68401 235989
rect 68429 235961 68464 235989
rect 68304 235944 68464 235961
rect 83664 236175 83824 236192
rect 83664 236147 83699 236175
rect 83727 236147 83761 236175
rect 83789 236147 83824 236175
rect 83664 236113 83824 236147
rect 83664 236085 83699 236113
rect 83727 236085 83761 236113
rect 83789 236085 83824 236113
rect 83664 236051 83824 236085
rect 83664 236023 83699 236051
rect 83727 236023 83761 236051
rect 83789 236023 83824 236051
rect 83664 235989 83824 236023
rect 83664 235961 83699 235989
rect 83727 235961 83761 235989
rect 83789 235961 83824 235989
rect 83664 235944 83824 235961
rect 94869 236175 95179 244961
rect 94869 236147 94917 236175
rect 94945 236147 94979 236175
rect 95007 236147 95041 236175
rect 95069 236147 95103 236175
rect 95131 236147 95179 236175
rect 94869 236113 95179 236147
rect 94869 236085 94917 236113
rect 94945 236085 94979 236113
rect 95007 236085 95041 236113
rect 95069 236085 95103 236113
rect 95131 236085 95179 236113
rect 94869 236051 95179 236085
rect 94869 236023 94917 236051
rect 94945 236023 94979 236051
rect 95007 236023 95041 236051
rect 95069 236023 95103 236051
rect 95131 236023 95179 236051
rect 94869 235989 95179 236023
rect 94869 235961 94917 235989
rect 94945 235961 94979 235989
rect 95007 235961 95041 235989
rect 95069 235961 95103 235989
rect 95131 235961 95179 235989
rect 29904 230175 30064 230192
rect 29904 230147 29939 230175
rect 29967 230147 30001 230175
rect 30029 230147 30064 230175
rect 29904 230113 30064 230147
rect 29904 230085 29939 230113
rect 29967 230085 30001 230113
rect 30029 230085 30064 230113
rect 29904 230051 30064 230085
rect 29904 230023 29939 230051
rect 29967 230023 30001 230051
rect 30029 230023 30064 230051
rect 29904 229989 30064 230023
rect 29904 229961 29939 229989
rect 29967 229961 30001 229989
rect 30029 229961 30064 229989
rect 29904 229944 30064 229961
rect 45264 230175 45424 230192
rect 45264 230147 45299 230175
rect 45327 230147 45361 230175
rect 45389 230147 45424 230175
rect 45264 230113 45424 230147
rect 45264 230085 45299 230113
rect 45327 230085 45361 230113
rect 45389 230085 45424 230113
rect 45264 230051 45424 230085
rect 45264 230023 45299 230051
rect 45327 230023 45361 230051
rect 45389 230023 45424 230051
rect 45264 229989 45424 230023
rect 45264 229961 45299 229989
rect 45327 229961 45361 229989
rect 45389 229961 45424 229989
rect 45264 229944 45424 229961
rect 60624 230175 60784 230192
rect 60624 230147 60659 230175
rect 60687 230147 60721 230175
rect 60749 230147 60784 230175
rect 60624 230113 60784 230147
rect 60624 230085 60659 230113
rect 60687 230085 60721 230113
rect 60749 230085 60784 230113
rect 60624 230051 60784 230085
rect 60624 230023 60659 230051
rect 60687 230023 60721 230051
rect 60749 230023 60784 230051
rect 60624 229989 60784 230023
rect 60624 229961 60659 229989
rect 60687 229961 60721 229989
rect 60749 229961 60784 229989
rect 60624 229944 60784 229961
rect 75984 230175 76144 230192
rect 75984 230147 76019 230175
rect 76047 230147 76081 230175
rect 76109 230147 76144 230175
rect 75984 230113 76144 230147
rect 75984 230085 76019 230113
rect 76047 230085 76081 230113
rect 76109 230085 76144 230113
rect 75984 230051 76144 230085
rect 75984 230023 76019 230051
rect 76047 230023 76081 230051
rect 76109 230023 76144 230051
rect 75984 229989 76144 230023
rect 75984 229961 76019 229989
rect 76047 229961 76081 229989
rect 76109 229961 76144 229989
rect 75984 229944 76144 229961
rect 18069 227147 18117 227175
rect 18145 227147 18179 227175
rect 18207 227147 18241 227175
rect 18269 227147 18303 227175
rect 18331 227147 18379 227175
rect 18069 227113 18379 227147
rect 18069 227085 18117 227113
rect 18145 227085 18179 227113
rect 18207 227085 18241 227113
rect 18269 227085 18303 227113
rect 18331 227085 18379 227113
rect 18069 227051 18379 227085
rect 18069 227023 18117 227051
rect 18145 227023 18179 227051
rect 18207 227023 18241 227051
rect 18269 227023 18303 227051
rect 18331 227023 18379 227051
rect 18069 226989 18379 227023
rect 18069 226961 18117 226989
rect 18145 226961 18179 226989
rect 18207 226961 18241 226989
rect 18269 226961 18303 226989
rect 18331 226961 18379 226989
rect 18069 218175 18379 226961
rect 22224 227175 22384 227192
rect 22224 227147 22259 227175
rect 22287 227147 22321 227175
rect 22349 227147 22384 227175
rect 22224 227113 22384 227147
rect 22224 227085 22259 227113
rect 22287 227085 22321 227113
rect 22349 227085 22384 227113
rect 22224 227051 22384 227085
rect 22224 227023 22259 227051
rect 22287 227023 22321 227051
rect 22349 227023 22384 227051
rect 22224 226989 22384 227023
rect 22224 226961 22259 226989
rect 22287 226961 22321 226989
rect 22349 226961 22384 226989
rect 22224 226944 22384 226961
rect 37584 227175 37744 227192
rect 37584 227147 37619 227175
rect 37647 227147 37681 227175
rect 37709 227147 37744 227175
rect 37584 227113 37744 227147
rect 37584 227085 37619 227113
rect 37647 227085 37681 227113
rect 37709 227085 37744 227113
rect 37584 227051 37744 227085
rect 37584 227023 37619 227051
rect 37647 227023 37681 227051
rect 37709 227023 37744 227051
rect 37584 226989 37744 227023
rect 37584 226961 37619 226989
rect 37647 226961 37681 226989
rect 37709 226961 37744 226989
rect 37584 226944 37744 226961
rect 52944 227175 53104 227192
rect 52944 227147 52979 227175
rect 53007 227147 53041 227175
rect 53069 227147 53104 227175
rect 52944 227113 53104 227147
rect 52944 227085 52979 227113
rect 53007 227085 53041 227113
rect 53069 227085 53104 227113
rect 52944 227051 53104 227085
rect 52944 227023 52979 227051
rect 53007 227023 53041 227051
rect 53069 227023 53104 227051
rect 52944 226989 53104 227023
rect 52944 226961 52979 226989
rect 53007 226961 53041 226989
rect 53069 226961 53104 226989
rect 52944 226944 53104 226961
rect 68304 227175 68464 227192
rect 68304 227147 68339 227175
rect 68367 227147 68401 227175
rect 68429 227147 68464 227175
rect 68304 227113 68464 227147
rect 68304 227085 68339 227113
rect 68367 227085 68401 227113
rect 68429 227085 68464 227113
rect 68304 227051 68464 227085
rect 68304 227023 68339 227051
rect 68367 227023 68401 227051
rect 68429 227023 68464 227051
rect 68304 226989 68464 227023
rect 68304 226961 68339 226989
rect 68367 226961 68401 226989
rect 68429 226961 68464 226989
rect 68304 226944 68464 226961
rect 83664 227175 83824 227192
rect 83664 227147 83699 227175
rect 83727 227147 83761 227175
rect 83789 227147 83824 227175
rect 83664 227113 83824 227147
rect 83664 227085 83699 227113
rect 83727 227085 83761 227113
rect 83789 227085 83824 227113
rect 83664 227051 83824 227085
rect 83664 227023 83699 227051
rect 83727 227023 83761 227051
rect 83789 227023 83824 227051
rect 83664 226989 83824 227023
rect 83664 226961 83699 226989
rect 83727 226961 83761 226989
rect 83789 226961 83824 226989
rect 83664 226944 83824 226961
rect 94869 227175 95179 235961
rect 94869 227147 94917 227175
rect 94945 227147 94979 227175
rect 95007 227147 95041 227175
rect 95069 227147 95103 227175
rect 95131 227147 95179 227175
rect 94869 227113 95179 227147
rect 94869 227085 94917 227113
rect 94945 227085 94979 227113
rect 95007 227085 95041 227113
rect 95069 227085 95103 227113
rect 95131 227085 95179 227113
rect 94869 227051 95179 227085
rect 94869 227023 94917 227051
rect 94945 227023 94979 227051
rect 95007 227023 95041 227051
rect 95069 227023 95103 227051
rect 95131 227023 95179 227051
rect 94869 226989 95179 227023
rect 94869 226961 94917 226989
rect 94945 226961 94979 226989
rect 95007 226961 95041 226989
rect 95069 226961 95103 226989
rect 95131 226961 95179 226989
rect 29904 221175 30064 221192
rect 29904 221147 29939 221175
rect 29967 221147 30001 221175
rect 30029 221147 30064 221175
rect 29904 221113 30064 221147
rect 29904 221085 29939 221113
rect 29967 221085 30001 221113
rect 30029 221085 30064 221113
rect 29904 221051 30064 221085
rect 29904 221023 29939 221051
rect 29967 221023 30001 221051
rect 30029 221023 30064 221051
rect 29904 220989 30064 221023
rect 29904 220961 29939 220989
rect 29967 220961 30001 220989
rect 30029 220961 30064 220989
rect 29904 220944 30064 220961
rect 45264 221175 45424 221192
rect 45264 221147 45299 221175
rect 45327 221147 45361 221175
rect 45389 221147 45424 221175
rect 45264 221113 45424 221147
rect 45264 221085 45299 221113
rect 45327 221085 45361 221113
rect 45389 221085 45424 221113
rect 45264 221051 45424 221085
rect 45264 221023 45299 221051
rect 45327 221023 45361 221051
rect 45389 221023 45424 221051
rect 45264 220989 45424 221023
rect 45264 220961 45299 220989
rect 45327 220961 45361 220989
rect 45389 220961 45424 220989
rect 45264 220944 45424 220961
rect 60624 221175 60784 221192
rect 60624 221147 60659 221175
rect 60687 221147 60721 221175
rect 60749 221147 60784 221175
rect 60624 221113 60784 221147
rect 60624 221085 60659 221113
rect 60687 221085 60721 221113
rect 60749 221085 60784 221113
rect 60624 221051 60784 221085
rect 60624 221023 60659 221051
rect 60687 221023 60721 221051
rect 60749 221023 60784 221051
rect 60624 220989 60784 221023
rect 60624 220961 60659 220989
rect 60687 220961 60721 220989
rect 60749 220961 60784 220989
rect 60624 220944 60784 220961
rect 75984 221175 76144 221192
rect 75984 221147 76019 221175
rect 76047 221147 76081 221175
rect 76109 221147 76144 221175
rect 75984 221113 76144 221147
rect 75984 221085 76019 221113
rect 76047 221085 76081 221113
rect 76109 221085 76144 221113
rect 75984 221051 76144 221085
rect 75984 221023 76019 221051
rect 76047 221023 76081 221051
rect 76109 221023 76144 221051
rect 75984 220989 76144 221023
rect 75984 220961 76019 220989
rect 76047 220961 76081 220989
rect 76109 220961 76144 220989
rect 75984 220944 76144 220961
rect 18069 218147 18117 218175
rect 18145 218147 18179 218175
rect 18207 218147 18241 218175
rect 18269 218147 18303 218175
rect 18331 218147 18379 218175
rect 18069 218113 18379 218147
rect 18069 218085 18117 218113
rect 18145 218085 18179 218113
rect 18207 218085 18241 218113
rect 18269 218085 18303 218113
rect 18331 218085 18379 218113
rect 18069 218051 18379 218085
rect 18069 218023 18117 218051
rect 18145 218023 18179 218051
rect 18207 218023 18241 218051
rect 18269 218023 18303 218051
rect 18331 218023 18379 218051
rect 18069 217989 18379 218023
rect 18069 217961 18117 217989
rect 18145 217961 18179 217989
rect 18207 217961 18241 217989
rect 18269 217961 18303 217989
rect 18331 217961 18379 217989
rect 5558 151601 5586 151606
rect 5614 215978 5642 215983
rect 5614 149954 5642 215950
rect 18069 209175 18379 217961
rect 22224 218175 22384 218192
rect 22224 218147 22259 218175
rect 22287 218147 22321 218175
rect 22349 218147 22384 218175
rect 22224 218113 22384 218147
rect 22224 218085 22259 218113
rect 22287 218085 22321 218113
rect 22349 218085 22384 218113
rect 22224 218051 22384 218085
rect 22224 218023 22259 218051
rect 22287 218023 22321 218051
rect 22349 218023 22384 218051
rect 22224 217989 22384 218023
rect 22224 217961 22259 217989
rect 22287 217961 22321 217989
rect 22349 217961 22384 217989
rect 22224 217944 22384 217961
rect 37584 218175 37744 218192
rect 37584 218147 37619 218175
rect 37647 218147 37681 218175
rect 37709 218147 37744 218175
rect 37584 218113 37744 218147
rect 37584 218085 37619 218113
rect 37647 218085 37681 218113
rect 37709 218085 37744 218113
rect 37584 218051 37744 218085
rect 37584 218023 37619 218051
rect 37647 218023 37681 218051
rect 37709 218023 37744 218051
rect 37584 217989 37744 218023
rect 37584 217961 37619 217989
rect 37647 217961 37681 217989
rect 37709 217961 37744 217989
rect 37584 217944 37744 217961
rect 52944 218175 53104 218192
rect 52944 218147 52979 218175
rect 53007 218147 53041 218175
rect 53069 218147 53104 218175
rect 52944 218113 53104 218147
rect 52944 218085 52979 218113
rect 53007 218085 53041 218113
rect 53069 218085 53104 218113
rect 52944 218051 53104 218085
rect 52944 218023 52979 218051
rect 53007 218023 53041 218051
rect 53069 218023 53104 218051
rect 52944 217989 53104 218023
rect 52944 217961 52979 217989
rect 53007 217961 53041 217989
rect 53069 217961 53104 217989
rect 52944 217944 53104 217961
rect 68304 218175 68464 218192
rect 68304 218147 68339 218175
rect 68367 218147 68401 218175
rect 68429 218147 68464 218175
rect 68304 218113 68464 218147
rect 68304 218085 68339 218113
rect 68367 218085 68401 218113
rect 68429 218085 68464 218113
rect 68304 218051 68464 218085
rect 68304 218023 68339 218051
rect 68367 218023 68401 218051
rect 68429 218023 68464 218051
rect 68304 217989 68464 218023
rect 68304 217961 68339 217989
rect 68367 217961 68401 217989
rect 68429 217961 68464 217989
rect 68304 217944 68464 217961
rect 83664 218175 83824 218192
rect 83664 218147 83699 218175
rect 83727 218147 83761 218175
rect 83789 218147 83824 218175
rect 83664 218113 83824 218147
rect 83664 218085 83699 218113
rect 83727 218085 83761 218113
rect 83789 218085 83824 218113
rect 83664 218051 83824 218085
rect 83664 218023 83699 218051
rect 83727 218023 83761 218051
rect 83789 218023 83824 218051
rect 83664 217989 83824 218023
rect 83664 217961 83699 217989
rect 83727 217961 83761 217989
rect 83789 217961 83824 217989
rect 83664 217944 83824 217961
rect 94869 218175 95179 226961
rect 94869 218147 94917 218175
rect 94945 218147 94979 218175
rect 95007 218147 95041 218175
rect 95069 218147 95103 218175
rect 95131 218147 95179 218175
rect 94869 218113 95179 218147
rect 94869 218085 94917 218113
rect 94945 218085 94979 218113
rect 95007 218085 95041 218113
rect 95069 218085 95103 218113
rect 95131 218085 95179 218113
rect 94869 218051 95179 218085
rect 94869 218023 94917 218051
rect 94945 218023 94979 218051
rect 95007 218023 95041 218051
rect 95069 218023 95103 218051
rect 95131 218023 95179 218051
rect 94869 217989 95179 218023
rect 94869 217961 94917 217989
rect 94945 217961 94979 217989
rect 95007 217961 95041 217989
rect 95069 217961 95103 217989
rect 95131 217961 95179 217989
rect 29904 212175 30064 212192
rect 29904 212147 29939 212175
rect 29967 212147 30001 212175
rect 30029 212147 30064 212175
rect 29904 212113 30064 212147
rect 29904 212085 29939 212113
rect 29967 212085 30001 212113
rect 30029 212085 30064 212113
rect 29904 212051 30064 212085
rect 29904 212023 29939 212051
rect 29967 212023 30001 212051
rect 30029 212023 30064 212051
rect 29904 211989 30064 212023
rect 29904 211961 29939 211989
rect 29967 211961 30001 211989
rect 30029 211961 30064 211989
rect 29904 211944 30064 211961
rect 45264 212175 45424 212192
rect 45264 212147 45299 212175
rect 45327 212147 45361 212175
rect 45389 212147 45424 212175
rect 45264 212113 45424 212147
rect 45264 212085 45299 212113
rect 45327 212085 45361 212113
rect 45389 212085 45424 212113
rect 45264 212051 45424 212085
rect 45264 212023 45299 212051
rect 45327 212023 45361 212051
rect 45389 212023 45424 212051
rect 45264 211989 45424 212023
rect 45264 211961 45299 211989
rect 45327 211961 45361 211989
rect 45389 211961 45424 211989
rect 45264 211944 45424 211961
rect 60624 212175 60784 212192
rect 60624 212147 60659 212175
rect 60687 212147 60721 212175
rect 60749 212147 60784 212175
rect 60624 212113 60784 212147
rect 60624 212085 60659 212113
rect 60687 212085 60721 212113
rect 60749 212085 60784 212113
rect 60624 212051 60784 212085
rect 60624 212023 60659 212051
rect 60687 212023 60721 212051
rect 60749 212023 60784 212051
rect 60624 211989 60784 212023
rect 60624 211961 60659 211989
rect 60687 211961 60721 211989
rect 60749 211961 60784 211989
rect 60624 211944 60784 211961
rect 75984 212175 76144 212192
rect 75984 212147 76019 212175
rect 76047 212147 76081 212175
rect 76109 212147 76144 212175
rect 75984 212113 76144 212147
rect 75984 212085 76019 212113
rect 76047 212085 76081 212113
rect 76109 212085 76144 212113
rect 75984 212051 76144 212085
rect 75984 212023 76019 212051
rect 76047 212023 76081 212051
rect 76109 212023 76144 212051
rect 75984 211989 76144 212023
rect 75984 211961 76019 211989
rect 76047 211961 76081 211989
rect 76109 211961 76144 211989
rect 75984 211944 76144 211961
rect 18069 209147 18117 209175
rect 18145 209147 18179 209175
rect 18207 209147 18241 209175
rect 18269 209147 18303 209175
rect 18331 209147 18379 209175
rect 18069 209113 18379 209147
rect 18069 209085 18117 209113
rect 18145 209085 18179 209113
rect 18207 209085 18241 209113
rect 18269 209085 18303 209113
rect 18331 209085 18379 209113
rect 18069 209051 18379 209085
rect 18069 209023 18117 209051
rect 18145 209023 18179 209051
rect 18207 209023 18241 209051
rect 18269 209023 18303 209051
rect 18331 209023 18379 209051
rect 18069 208989 18379 209023
rect 18069 208961 18117 208989
rect 18145 208961 18179 208989
rect 18207 208961 18241 208989
rect 18269 208961 18303 208989
rect 18331 208961 18379 208989
rect 5614 149921 5642 149926
rect 6286 201866 6314 201871
rect 6286 148834 6314 201838
rect 18069 200175 18379 208961
rect 22224 209175 22384 209192
rect 22224 209147 22259 209175
rect 22287 209147 22321 209175
rect 22349 209147 22384 209175
rect 22224 209113 22384 209147
rect 22224 209085 22259 209113
rect 22287 209085 22321 209113
rect 22349 209085 22384 209113
rect 22224 209051 22384 209085
rect 22224 209023 22259 209051
rect 22287 209023 22321 209051
rect 22349 209023 22384 209051
rect 22224 208989 22384 209023
rect 22224 208961 22259 208989
rect 22287 208961 22321 208989
rect 22349 208961 22384 208989
rect 22224 208944 22384 208961
rect 37584 209175 37744 209192
rect 37584 209147 37619 209175
rect 37647 209147 37681 209175
rect 37709 209147 37744 209175
rect 37584 209113 37744 209147
rect 37584 209085 37619 209113
rect 37647 209085 37681 209113
rect 37709 209085 37744 209113
rect 37584 209051 37744 209085
rect 37584 209023 37619 209051
rect 37647 209023 37681 209051
rect 37709 209023 37744 209051
rect 37584 208989 37744 209023
rect 37584 208961 37619 208989
rect 37647 208961 37681 208989
rect 37709 208961 37744 208989
rect 37584 208944 37744 208961
rect 52944 209175 53104 209192
rect 52944 209147 52979 209175
rect 53007 209147 53041 209175
rect 53069 209147 53104 209175
rect 52944 209113 53104 209147
rect 52944 209085 52979 209113
rect 53007 209085 53041 209113
rect 53069 209085 53104 209113
rect 52944 209051 53104 209085
rect 52944 209023 52979 209051
rect 53007 209023 53041 209051
rect 53069 209023 53104 209051
rect 52944 208989 53104 209023
rect 52944 208961 52979 208989
rect 53007 208961 53041 208989
rect 53069 208961 53104 208989
rect 52944 208944 53104 208961
rect 68304 209175 68464 209192
rect 68304 209147 68339 209175
rect 68367 209147 68401 209175
rect 68429 209147 68464 209175
rect 68304 209113 68464 209147
rect 68304 209085 68339 209113
rect 68367 209085 68401 209113
rect 68429 209085 68464 209113
rect 68304 209051 68464 209085
rect 68304 209023 68339 209051
rect 68367 209023 68401 209051
rect 68429 209023 68464 209051
rect 68304 208989 68464 209023
rect 68304 208961 68339 208989
rect 68367 208961 68401 208989
rect 68429 208961 68464 208989
rect 68304 208944 68464 208961
rect 83664 209175 83824 209192
rect 83664 209147 83699 209175
rect 83727 209147 83761 209175
rect 83789 209147 83824 209175
rect 83664 209113 83824 209147
rect 83664 209085 83699 209113
rect 83727 209085 83761 209113
rect 83789 209085 83824 209113
rect 83664 209051 83824 209085
rect 83664 209023 83699 209051
rect 83727 209023 83761 209051
rect 83789 209023 83824 209051
rect 83664 208989 83824 209023
rect 83664 208961 83699 208989
rect 83727 208961 83761 208989
rect 83789 208961 83824 208989
rect 83664 208944 83824 208961
rect 94869 209175 95179 217961
rect 94869 209147 94917 209175
rect 94945 209147 94979 209175
rect 95007 209147 95041 209175
rect 95069 209147 95103 209175
rect 95131 209147 95179 209175
rect 94869 209113 95179 209147
rect 94869 209085 94917 209113
rect 94945 209085 94979 209113
rect 95007 209085 95041 209113
rect 95069 209085 95103 209113
rect 95131 209085 95179 209113
rect 94869 209051 95179 209085
rect 94869 209023 94917 209051
rect 94945 209023 94979 209051
rect 95007 209023 95041 209051
rect 95069 209023 95103 209051
rect 95131 209023 95179 209051
rect 94869 208989 95179 209023
rect 94869 208961 94917 208989
rect 94945 208961 94979 208989
rect 95007 208961 95041 208989
rect 95069 208961 95103 208989
rect 95131 208961 95179 208989
rect 29904 203175 30064 203192
rect 29904 203147 29939 203175
rect 29967 203147 30001 203175
rect 30029 203147 30064 203175
rect 29904 203113 30064 203147
rect 29904 203085 29939 203113
rect 29967 203085 30001 203113
rect 30029 203085 30064 203113
rect 29904 203051 30064 203085
rect 29904 203023 29939 203051
rect 29967 203023 30001 203051
rect 30029 203023 30064 203051
rect 29904 202989 30064 203023
rect 29904 202961 29939 202989
rect 29967 202961 30001 202989
rect 30029 202961 30064 202989
rect 29904 202944 30064 202961
rect 45264 203175 45424 203192
rect 45264 203147 45299 203175
rect 45327 203147 45361 203175
rect 45389 203147 45424 203175
rect 45264 203113 45424 203147
rect 45264 203085 45299 203113
rect 45327 203085 45361 203113
rect 45389 203085 45424 203113
rect 45264 203051 45424 203085
rect 45264 203023 45299 203051
rect 45327 203023 45361 203051
rect 45389 203023 45424 203051
rect 45264 202989 45424 203023
rect 45264 202961 45299 202989
rect 45327 202961 45361 202989
rect 45389 202961 45424 202989
rect 45264 202944 45424 202961
rect 60624 203175 60784 203192
rect 60624 203147 60659 203175
rect 60687 203147 60721 203175
rect 60749 203147 60784 203175
rect 60624 203113 60784 203147
rect 60624 203085 60659 203113
rect 60687 203085 60721 203113
rect 60749 203085 60784 203113
rect 60624 203051 60784 203085
rect 60624 203023 60659 203051
rect 60687 203023 60721 203051
rect 60749 203023 60784 203051
rect 60624 202989 60784 203023
rect 60624 202961 60659 202989
rect 60687 202961 60721 202989
rect 60749 202961 60784 202989
rect 60624 202944 60784 202961
rect 75984 203175 76144 203192
rect 75984 203147 76019 203175
rect 76047 203147 76081 203175
rect 76109 203147 76144 203175
rect 75984 203113 76144 203147
rect 75984 203085 76019 203113
rect 76047 203085 76081 203113
rect 76109 203085 76144 203113
rect 75984 203051 76144 203085
rect 75984 203023 76019 203051
rect 76047 203023 76081 203051
rect 76109 203023 76144 203051
rect 75984 202989 76144 203023
rect 75984 202961 76019 202989
rect 76047 202961 76081 202989
rect 76109 202961 76144 202989
rect 75984 202944 76144 202961
rect 18069 200147 18117 200175
rect 18145 200147 18179 200175
rect 18207 200147 18241 200175
rect 18269 200147 18303 200175
rect 18331 200147 18379 200175
rect 18069 200113 18379 200147
rect 18069 200085 18117 200113
rect 18145 200085 18179 200113
rect 18207 200085 18241 200113
rect 18269 200085 18303 200113
rect 18331 200085 18379 200113
rect 18069 200051 18379 200085
rect 18069 200023 18117 200051
rect 18145 200023 18179 200051
rect 18207 200023 18241 200051
rect 18269 200023 18303 200051
rect 18331 200023 18379 200051
rect 18069 199989 18379 200023
rect 18069 199961 18117 199989
rect 18145 199961 18179 199989
rect 18207 199961 18241 199989
rect 18269 199961 18303 199989
rect 18331 199961 18379 199989
rect 6286 148801 6314 148806
rect 6342 194810 6370 194815
rect 6342 148274 6370 194782
rect 18069 191175 18379 199961
rect 22224 200175 22384 200192
rect 22224 200147 22259 200175
rect 22287 200147 22321 200175
rect 22349 200147 22384 200175
rect 22224 200113 22384 200147
rect 22224 200085 22259 200113
rect 22287 200085 22321 200113
rect 22349 200085 22384 200113
rect 22224 200051 22384 200085
rect 22224 200023 22259 200051
rect 22287 200023 22321 200051
rect 22349 200023 22384 200051
rect 22224 199989 22384 200023
rect 22224 199961 22259 199989
rect 22287 199961 22321 199989
rect 22349 199961 22384 199989
rect 22224 199944 22384 199961
rect 37584 200175 37744 200192
rect 37584 200147 37619 200175
rect 37647 200147 37681 200175
rect 37709 200147 37744 200175
rect 37584 200113 37744 200147
rect 37584 200085 37619 200113
rect 37647 200085 37681 200113
rect 37709 200085 37744 200113
rect 37584 200051 37744 200085
rect 37584 200023 37619 200051
rect 37647 200023 37681 200051
rect 37709 200023 37744 200051
rect 37584 199989 37744 200023
rect 37584 199961 37619 199989
rect 37647 199961 37681 199989
rect 37709 199961 37744 199989
rect 37584 199944 37744 199961
rect 52944 200175 53104 200192
rect 52944 200147 52979 200175
rect 53007 200147 53041 200175
rect 53069 200147 53104 200175
rect 52944 200113 53104 200147
rect 52944 200085 52979 200113
rect 53007 200085 53041 200113
rect 53069 200085 53104 200113
rect 52944 200051 53104 200085
rect 52944 200023 52979 200051
rect 53007 200023 53041 200051
rect 53069 200023 53104 200051
rect 52944 199989 53104 200023
rect 52944 199961 52979 199989
rect 53007 199961 53041 199989
rect 53069 199961 53104 199989
rect 52944 199944 53104 199961
rect 68304 200175 68464 200192
rect 68304 200147 68339 200175
rect 68367 200147 68401 200175
rect 68429 200147 68464 200175
rect 68304 200113 68464 200147
rect 68304 200085 68339 200113
rect 68367 200085 68401 200113
rect 68429 200085 68464 200113
rect 68304 200051 68464 200085
rect 68304 200023 68339 200051
rect 68367 200023 68401 200051
rect 68429 200023 68464 200051
rect 68304 199989 68464 200023
rect 68304 199961 68339 199989
rect 68367 199961 68401 199989
rect 68429 199961 68464 199989
rect 68304 199944 68464 199961
rect 83664 200175 83824 200192
rect 83664 200147 83699 200175
rect 83727 200147 83761 200175
rect 83789 200147 83824 200175
rect 83664 200113 83824 200147
rect 83664 200085 83699 200113
rect 83727 200085 83761 200113
rect 83789 200085 83824 200113
rect 83664 200051 83824 200085
rect 83664 200023 83699 200051
rect 83727 200023 83761 200051
rect 83789 200023 83824 200051
rect 83664 199989 83824 200023
rect 83664 199961 83699 199989
rect 83727 199961 83761 199989
rect 83789 199961 83824 199989
rect 83664 199944 83824 199961
rect 94869 200175 95179 208961
rect 94869 200147 94917 200175
rect 94945 200147 94979 200175
rect 95007 200147 95041 200175
rect 95069 200147 95103 200175
rect 95131 200147 95179 200175
rect 94869 200113 95179 200147
rect 94869 200085 94917 200113
rect 94945 200085 94979 200113
rect 95007 200085 95041 200113
rect 95069 200085 95103 200113
rect 95131 200085 95179 200113
rect 94869 200051 95179 200085
rect 94869 200023 94917 200051
rect 94945 200023 94979 200051
rect 95007 200023 95041 200051
rect 95069 200023 95103 200051
rect 95131 200023 95179 200051
rect 94869 199989 95179 200023
rect 94869 199961 94917 199989
rect 94945 199961 94979 199989
rect 95007 199961 95041 199989
rect 95069 199961 95103 199989
rect 95131 199961 95179 199989
rect 29904 194175 30064 194192
rect 29904 194147 29939 194175
rect 29967 194147 30001 194175
rect 30029 194147 30064 194175
rect 29904 194113 30064 194147
rect 29904 194085 29939 194113
rect 29967 194085 30001 194113
rect 30029 194085 30064 194113
rect 29904 194051 30064 194085
rect 29904 194023 29939 194051
rect 29967 194023 30001 194051
rect 30029 194023 30064 194051
rect 29904 193989 30064 194023
rect 29904 193961 29939 193989
rect 29967 193961 30001 193989
rect 30029 193961 30064 193989
rect 29904 193944 30064 193961
rect 45264 194175 45424 194192
rect 45264 194147 45299 194175
rect 45327 194147 45361 194175
rect 45389 194147 45424 194175
rect 45264 194113 45424 194147
rect 45264 194085 45299 194113
rect 45327 194085 45361 194113
rect 45389 194085 45424 194113
rect 45264 194051 45424 194085
rect 45264 194023 45299 194051
rect 45327 194023 45361 194051
rect 45389 194023 45424 194051
rect 45264 193989 45424 194023
rect 45264 193961 45299 193989
rect 45327 193961 45361 193989
rect 45389 193961 45424 193989
rect 45264 193944 45424 193961
rect 60624 194175 60784 194192
rect 60624 194147 60659 194175
rect 60687 194147 60721 194175
rect 60749 194147 60784 194175
rect 60624 194113 60784 194147
rect 60624 194085 60659 194113
rect 60687 194085 60721 194113
rect 60749 194085 60784 194113
rect 60624 194051 60784 194085
rect 60624 194023 60659 194051
rect 60687 194023 60721 194051
rect 60749 194023 60784 194051
rect 60624 193989 60784 194023
rect 60624 193961 60659 193989
rect 60687 193961 60721 193989
rect 60749 193961 60784 193989
rect 60624 193944 60784 193961
rect 75984 194175 76144 194192
rect 75984 194147 76019 194175
rect 76047 194147 76081 194175
rect 76109 194147 76144 194175
rect 75984 194113 76144 194147
rect 75984 194085 76019 194113
rect 76047 194085 76081 194113
rect 76109 194085 76144 194113
rect 75984 194051 76144 194085
rect 75984 194023 76019 194051
rect 76047 194023 76081 194051
rect 76109 194023 76144 194051
rect 75984 193989 76144 194023
rect 75984 193961 76019 193989
rect 76047 193961 76081 193989
rect 76109 193961 76144 193989
rect 75984 193944 76144 193961
rect 18069 191147 18117 191175
rect 18145 191147 18179 191175
rect 18207 191147 18241 191175
rect 18269 191147 18303 191175
rect 18331 191147 18379 191175
rect 18069 191113 18379 191147
rect 18069 191085 18117 191113
rect 18145 191085 18179 191113
rect 18207 191085 18241 191113
rect 18269 191085 18303 191113
rect 18331 191085 18379 191113
rect 18069 191051 18379 191085
rect 18069 191023 18117 191051
rect 18145 191023 18179 191051
rect 18207 191023 18241 191051
rect 18269 191023 18303 191051
rect 18331 191023 18379 191051
rect 18069 190989 18379 191023
rect 18069 190961 18117 190989
rect 18145 190961 18179 190989
rect 18207 190961 18241 190989
rect 18269 190961 18303 190989
rect 18331 190961 18379 190989
rect 18069 182175 18379 190961
rect 22224 191175 22384 191192
rect 22224 191147 22259 191175
rect 22287 191147 22321 191175
rect 22349 191147 22384 191175
rect 22224 191113 22384 191147
rect 22224 191085 22259 191113
rect 22287 191085 22321 191113
rect 22349 191085 22384 191113
rect 22224 191051 22384 191085
rect 22224 191023 22259 191051
rect 22287 191023 22321 191051
rect 22349 191023 22384 191051
rect 22224 190989 22384 191023
rect 22224 190961 22259 190989
rect 22287 190961 22321 190989
rect 22349 190961 22384 190989
rect 22224 190944 22384 190961
rect 37584 191175 37744 191192
rect 37584 191147 37619 191175
rect 37647 191147 37681 191175
rect 37709 191147 37744 191175
rect 37584 191113 37744 191147
rect 37584 191085 37619 191113
rect 37647 191085 37681 191113
rect 37709 191085 37744 191113
rect 37584 191051 37744 191085
rect 37584 191023 37619 191051
rect 37647 191023 37681 191051
rect 37709 191023 37744 191051
rect 37584 190989 37744 191023
rect 37584 190961 37619 190989
rect 37647 190961 37681 190989
rect 37709 190961 37744 190989
rect 37584 190944 37744 190961
rect 52944 191175 53104 191192
rect 52944 191147 52979 191175
rect 53007 191147 53041 191175
rect 53069 191147 53104 191175
rect 52944 191113 53104 191147
rect 52944 191085 52979 191113
rect 53007 191085 53041 191113
rect 53069 191085 53104 191113
rect 52944 191051 53104 191085
rect 52944 191023 52979 191051
rect 53007 191023 53041 191051
rect 53069 191023 53104 191051
rect 52944 190989 53104 191023
rect 52944 190961 52979 190989
rect 53007 190961 53041 190989
rect 53069 190961 53104 190989
rect 52944 190944 53104 190961
rect 68304 191175 68464 191192
rect 68304 191147 68339 191175
rect 68367 191147 68401 191175
rect 68429 191147 68464 191175
rect 68304 191113 68464 191147
rect 68304 191085 68339 191113
rect 68367 191085 68401 191113
rect 68429 191085 68464 191113
rect 68304 191051 68464 191085
rect 68304 191023 68339 191051
rect 68367 191023 68401 191051
rect 68429 191023 68464 191051
rect 68304 190989 68464 191023
rect 68304 190961 68339 190989
rect 68367 190961 68401 190989
rect 68429 190961 68464 190989
rect 68304 190944 68464 190961
rect 83664 191175 83824 191192
rect 83664 191147 83699 191175
rect 83727 191147 83761 191175
rect 83789 191147 83824 191175
rect 83664 191113 83824 191147
rect 83664 191085 83699 191113
rect 83727 191085 83761 191113
rect 83789 191085 83824 191113
rect 83664 191051 83824 191085
rect 83664 191023 83699 191051
rect 83727 191023 83761 191051
rect 83789 191023 83824 191051
rect 83664 190989 83824 191023
rect 83664 190961 83699 190989
rect 83727 190961 83761 190989
rect 83789 190961 83824 190989
rect 83664 190944 83824 190961
rect 94869 191175 95179 199961
rect 94869 191147 94917 191175
rect 94945 191147 94979 191175
rect 95007 191147 95041 191175
rect 95069 191147 95103 191175
rect 95131 191147 95179 191175
rect 94869 191113 95179 191147
rect 94869 191085 94917 191113
rect 94945 191085 94979 191113
rect 95007 191085 95041 191113
rect 95069 191085 95103 191113
rect 95131 191085 95179 191113
rect 94869 191051 95179 191085
rect 94869 191023 94917 191051
rect 94945 191023 94979 191051
rect 95007 191023 95041 191051
rect 95069 191023 95103 191051
rect 95131 191023 95179 191051
rect 94869 190989 95179 191023
rect 94869 190961 94917 190989
rect 94945 190961 94979 190989
rect 95007 190961 95041 190989
rect 95069 190961 95103 190989
rect 95131 190961 95179 190989
rect 29904 185175 30064 185192
rect 29904 185147 29939 185175
rect 29967 185147 30001 185175
rect 30029 185147 30064 185175
rect 29904 185113 30064 185147
rect 29904 185085 29939 185113
rect 29967 185085 30001 185113
rect 30029 185085 30064 185113
rect 29904 185051 30064 185085
rect 29904 185023 29939 185051
rect 29967 185023 30001 185051
rect 30029 185023 30064 185051
rect 29904 184989 30064 185023
rect 29904 184961 29939 184989
rect 29967 184961 30001 184989
rect 30029 184961 30064 184989
rect 29904 184944 30064 184961
rect 45264 185175 45424 185192
rect 45264 185147 45299 185175
rect 45327 185147 45361 185175
rect 45389 185147 45424 185175
rect 45264 185113 45424 185147
rect 45264 185085 45299 185113
rect 45327 185085 45361 185113
rect 45389 185085 45424 185113
rect 45264 185051 45424 185085
rect 45264 185023 45299 185051
rect 45327 185023 45361 185051
rect 45389 185023 45424 185051
rect 45264 184989 45424 185023
rect 45264 184961 45299 184989
rect 45327 184961 45361 184989
rect 45389 184961 45424 184989
rect 45264 184944 45424 184961
rect 60624 185175 60784 185192
rect 60624 185147 60659 185175
rect 60687 185147 60721 185175
rect 60749 185147 60784 185175
rect 60624 185113 60784 185147
rect 60624 185085 60659 185113
rect 60687 185085 60721 185113
rect 60749 185085 60784 185113
rect 60624 185051 60784 185085
rect 60624 185023 60659 185051
rect 60687 185023 60721 185051
rect 60749 185023 60784 185051
rect 60624 184989 60784 185023
rect 60624 184961 60659 184989
rect 60687 184961 60721 184989
rect 60749 184961 60784 184989
rect 60624 184944 60784 184961
rect 75984 185175 76144 185192
rect 75984 185147 76019 185175
rect 76047 185147 76081 185175
rect 76109 185147 76144 185175
rect 75984 185113 76144 185147
rect 75984 185085 76019 185113
rect 76047 185085 76081 185113
rect 76109 185085 76144 185113
rect 75984 185051 76144 185085
rect 75984 185023 76019 185051
rect 76047 185023 76081 185051
rect 76109 185023 76144 185051
rect 75984 184989 76144 185023
rect 75984 184961 76019 184989
rect 76047 184961 76081 184989
rect 76109 184961 76144 184989
rect 75984 184944 76144 184961
rect 18069 182147 18117 182175
rect 18145 182147 18179 182175
rect 18207 182147 18241 182175
rect 18269 182147 18303 182175
rect 18331 182147 18379 182175
rect 18069 182113 18379 182147
rect 18069 182085 18117 182113
rect 18145 182085 18179 182113
rect 18207 182085 18241 182113
rect 18269 182085 18303 182113
rect 18331 182085 18379 182113
rect 18069 182051 18379 182085
rect 18069 182023 18117 182051
rect 18145 182023 18179 182051
rect 18207 182023 18241 182051
rect 18269 182023 18303 182051
rect 18331 182023 18379 182051
rect 18069 181989 18379 182023
rect 18069 181961 18117 181989
rect 18145 181961 18179 181989
rect 18207 181961 18241 181989
rect 18269 181961 18303 181989
rect 18331 181961 18379 181989
rect 18069 173175 18379 181961
rect 22224 182175 22384 182192
rect 22224 182147 22259 182175
rect 22287 182147 22321 182175
rect 22349 182147 22384 182175
rect 22224 182113 22384 182147
rect 22224 182085 22259 182113
rect 22287 182085 22321 182113
rect 22349 182085 22384 182113
rect 22224 182051 22384 182085
rect 22224 182023 22259 182051
rect 22287 182023 22321 182051
rect 22349 182023 22384 182051
rect 22224 181989 22384 182023
rect 22224 181961 22259 181989
rect 22287 181961 22321 181989
rect 22349 181961 22384 181989
rect 22224 181944 22384 181961
rect 37584 182175 37744 182192
rect 37584 182147 37619 182175
rect 37647 182147 37681 182175
rect 37709 182147 37744 182175
rect 37584 182113 37744 182147
rect 37584 182085 37619 182113
rect 37647 182085 37681 182113
rect 37709 182085 37744 182113
rect 37584 182051 37744 182085
rect 37584 182023 37619 182051
rect 37647 182023 37681 182051
rect 37709 182023 37744 182051
rect 37584 181989 37744 182023
rect 37584 181961 37619 181989
rect 37647 181961 37681 181989
rect 37709 181961 37744 181989
rect 37584 181944 37744 181961
rect 52944 182175 53104 182192
rect 52944 182147 52979 182175
rect 53007 182147 53041 182175
rect 53069 182147 53104 182175
rect 52944 182113 53104 182147
rect 52944 182085 52979 182113
rect 53007 182085 53041 182113
rect 53069 182085 53104 182113
rect 52944 182051 53104 182085
rect 52944 182023 52979 182051
rect 53007 182023 53041 182051
rect 53069 182023 53104 182051
rect 52944 181989 53104 182023
rect 52944 181961 52979 181989
rect 53007 181961 53041 181989
rect 53069 181961 53104 181989
rect 52944 181944 53104 181961
rect 68304 182175 68464 182192
rect 68304 182147 68339 182175
rect 68367 182147 68401 182175
rect 68429 182147 68464 182175
rect 68304 182113 68464 182147
rect 68304 182085 68339 182113
rect 68367 182085 68401 182113
rect 68429 182085 68464 182113
rect 68304 182051 68464 182085
rect 68304 182023 68339 182051
rect 68367 182023 68401 182051
rect 68429 182023 68464 182051
rect 68304 181989 68464 182023
rect 68304 181961 68339 181989
rect 68367 181961 68401 181989
rect 68429 181961 68464 181989
rect 68304 181944 68464 181961
rect 83664 182175 83824 182192
rect 83664 182147 83699 182175
rect 83727 182147 83761 182175
rect 83789 182147 83824 182175
rect 83664 182113 83824 182147
rect 83664 182085 83699 182113
rect 83727 182085 83761 182113
rect 83789 182085 83824 182113
rect 83664 182051 83824 182085
rect 83664 182023 83699 182051
rect 83727 182023 83761 182051
rect 83789 182023 83824 182051
rect 83664 181989 83824 182023
rect 83664 181961 83699 181989
rect 83727 181961 83761 181989
rect 83789 181961 83824 181989
rect 83664 181944 83824 181961
rect 94869 182175 95179 190961
rect 94869 182147 94917 182175
rect 94945 182147 94979 182175
rect 95007 182147 95041 182175
rect 95069 182147 95103 182175
rect 95131 182147 95179 182175
rect 94869 182113 95179 182147
rect 94869 182085 94917 182113
rect 94945 182085 94979 182113
rect 95007 182085 95041 182113
rect 95069 182085 95103 182113
rect 95131 182085 95179 182113
rect 94869 182051 95179 182085
rect 94869 182023 94917 182051
rect 94945 182023 94979 182051
rect 95007 182023 95041 182051
rect 95069 182023 95103 182051
rect 95131 182023 95179 182051
rect 94869 181989 95179 182023
rect 94869 181961 94917 181989
rect 94945 181961 94979 181989
rect 95007 181961 95041 181989
rect 95069 181961 95103 181989
rect 95131 181961 95179 181989
rect 29904 176175 30064 176192
rect 29904 176147 29939 176175
rect 29967 176147 30001 176175
rect 30029 176147 30064 176175
rect 29904 176113 30064 176147
rect 29904 176085 29939 176113
rect 29967 176085 30001 176113
rect 30029 176085 30064 176113
rect 29904 176051 30064 176085
rect 29904 176023 29939 176051
rect 29967 176023 30001 176051
rect 30029 176023 30064 176051
rect 29904 175989 30064 176023
rect 29904 175961 29939 175989
rect 29967 175961 30001 175989
rect 30029 175961 30064 175989
rect 29904 175944 30064 175961
rect 45264 176175 45424 176192
rect 45264 176147 45299 176175
rect 45327 176147 45361 176175
rect 45389 176147 45424 176175
rect 45264 176113 45424 176147
rect 45264 176085 45299 176113
rect 45327 176085 45361 176113
rect 45389 176085 45424 176113
rect 45264 176051 45424 176085
rect 45264 176023 45299 176051
rect 45327 176023 45361 176051
rect 45389 176023 45424 176051
rect 45264 175989 45424 176023
rect 45264 175961 45299 175989
rect 45327 175961 45361 175989
rect 45389 175961 45424 175989
rect 45264 175944 45424 175961
rect 60624 176175 60784 176192
rect 60624 176147 60659 176175
rect 60687 176147 60721 176175
rect 60749 176147 60784 176175
rect 60624 176113 60784 176147
rect 60624 176085 60659 176113
rect 60687 176085 60721 176113
rect 60749 176085 60784 176113
rect 60624 176051 60784 176085
rect 60624 176023 60659 176051
rect 60687 176023 60721 176051
rect 60749 176023 60784 176051
rect 60624 175989 60784 176023
rect 60624 175961 60659 175989
rect 60687 175961 60721 175989
rect 60749 175961 60784 175989
rect 60624 175944 60784 175961
rect 75984 176175 76144 176192
rect 75984 176147 76019 176175
rect 76047 176147 76081 176175
rect 76109 176147 76144 176175
rect 75984 176113 76144 176147
rect 75984 176085 76019 176113
rect 76047 176085 76081 176113
rect 76109 176085 76144 176113
rect 75984 176051 76144 176085
rect 75984 176023 76019 176051
rect 76047 176023 76081 176051
rect 76109 176023 76144 176051
rect 75984 175989 76144 176023
rect 75984 175961 76019 175989
rect 76047 175961 76081 175989
rect 76109 175961 76144 175989
rect 75984 175944 76144 175961
rect 18069 173147 18117 173175
rect 18145 173147 18179 173175
rect 18207 173147 18241 173175
rect 18269 173147 18303 173175
rect 18331 173147 18379 173175
rect 18069 173113 18379 173147
rect 18069 173085 18117 173113
rect 18145 173085 18179 173113
rect 18207 173085 18241 173113
rect 18269 173085 18303 173113
rect 18331 173085 18379 173113
rect 18069 173051 18379 173085
rect 18069 173023 18117 173051
rect 18145 173023 18179 173051
rect 18207 173023 18241 173051
rect 18269 173023 18303 173051
rect 18331 173023 18379 173051
rect 18069 172989 18379 173023
rect 18069 172961 18117 172989
rect 18145 172961 18179 172989
rect 18207 172961 18241 172989
rect 18269 172961 18303 172989
rect 18331 172961 18379 172989
rect 18069 164175 18379 172961
rect 22224 173175 22384 173192
rect 22224 173147 22259 173175
rect 22287 173147 22321 173175
rect 22349 173147 22384 173175
rect 22224 173113 22384 173147
rect 22224 173085 22259 173113
rect 22287 173085 22321 173113
rect 22349 173085 22384 173113
rect 22224 173051 22384 173085
rect 22224 173023 22259 173051
rect 22287 173023 22321 173051
rect 22349 173023 22384 173051
rect 22224 172989 22384 173023
rect 22224 172961 22259 172989
rect 22287 172961 22321 172989
rect 22349 172961 22384 172989
rect 22224 172944 22384 172961
rect 37584 173175 37744 173192
rect 37584 173147 37619 173175
rect 37647 173147 37681 173175
rect 37709 173147 37744 173175
rect 37584 173113 37744 173147
rect 37584 173085 37619 173113
rect 37647 173085 37681 173113
rect 37709 173085 37744 173113
rect 37584 173051 37744 173085
rect 37584 173023 37619 173051
rect 37647 173023 37681 173051
rect 37709 173023 37744 173051
rect 37584 172989 37744 173023
rect 37584 172961 37619 172989
rect 37647 172961 37681 172989
rect 37709 172961 37744 172989
rect 37584 172944 37744 172961
rect 52944 173175 53104 173192
rect 52944 173147 52979 173175
rect 53007 173147 53041 173175
rect 53069 173147 53104 173175
rect 52944 173113 53104 173147
rect 52944 173085 52979 173113
rect 53007 173085 53041 173113
rect 53069 173085 53104 173113
rect 52944 173051 53104 173085
rect 52944 173023 52979 173051
rect 53007 173023 53041 173051
rect 53069 173023 53104 173051
rect 52944 172989 53104 173023
rect 52944 172961 52979 172989
rect 53007 172961 53041 172989
rect 53069 172961 53104 172989
rect 52944 172944 53104 172961
rect 68304 173175 68464 173192
rect 68304 173147 68339 173175
rect 68367 173147 68401 173175
rect 68429 173147 68464 173175
rect 68304 173113 68464 173147
rect 68304 173085 68339 173113
rect 68367 173085 68401 173113
rect 68429 173085 68464 173113
rect 68304 173051 68464 173085
rect 68304 173023 68339 173051
rect 68367 173023 68401 173051
rect 68429 173023 68464 173051
rect 68304 172989 68464 173023
rect 68304 172961 68339 172989
rect 68367 172961 68401 172989
rect 68429 172961 68464 172989
rect 68304 172944 68464 172961
rect 83664 173175 83824 173192
rect 83664 173147 83699 173175
rect 83727 173147 83761 173175
rect 83789 173147 83824 173175
rect 83664 173113 83824 173147
rect 83664 173085 83699 173113
rect 83727 173085 83761 173113
rect 83789 173085 83824 173113
rect 83664 173051 83824 173085
rect 83664 173023 83699 173051
rect 83727 173023 83761 173051
rect 83789 173023 83824 173051
rect 83664 172989 83824 173023
rect 83664 172961 83699 172989
rect 83727 172961 83761 172989
rect 83789 172961 83824 172989
rect 83664 172944 83824 172961
rect 94869 173175 95179 181961
rect 94869 173147 94917 173175
rect 94945 173147 94979 173175
rect 95007 173147 95041 173175
rect 95069 173147 95103 173175
rect 95131 173147 95179 173175
rect 94869 173113 95179 173147
rect 94869 173085 94917 173113
rect 94945 173085 94979 173113
rect 95007 173085 95041 173113
rect 95069 173085 95103 173113
rect 95131 173085 95179 173113
rect 94869 173051 95179 173085
rect 94869 173023 94917 173051
rect 94945 173023 94979 173051
rect 95007 173023 95041 173051
rect 95069 173023 95103 173051
rect 95131 173023 95179 173051
rect 94869 172989 95179 173023
rect 94869 172961 94917 172989
rect 94945 172961 94979 172989
rect 95007 172961 95041 172989
rect 95069 172961 95103 172989
rect 95131 172961 95179 172989
rect 18069 164147 18117 164175
rect 18145 164147 18179 164175
rect 18207 164147 18241 164175
rect 18269 164147 18303 164175
rect 18331 164147 18379 164175
rect 18069 164113 18379 164147
rect 18069 164085 18117 164113
rect 18145 164085 18179 164113
rect 18207 164085 18241 164113
rect 18269 164085 18303 164113
rect 18331 164085 18379 164113
rect 18069 164051 18379 164085
rect 18069 164023 18117 164051
rect 18145 164023 18179 164051
rect 18207 164023 18241 164051
rect 18269 164023 18303 164051
rect 18331 164023 18379 164051
rect 18069 163989 18379 164023
rect 18069 163961 18117 163989
rect 18145 163961 18179 163989
rect 18207 163961 18241 163989
rect 18269 163961 18303 163989
rect 18331 163961 18379 163989
rect 6342 148241 6370 148246
rect 6398 159530 6426 159535
rect 4942 147681 4970 147686
rect 6398 145474 6426 159502
rect 6398 145441 6426 145446
rect 18069 155175 18379 163961
rect 18069 155147 18117 155175
rect 18145 155147 18179 155175
rect 18207 155147 18241 155175
rect 18269 155147 18303 155175
rect 18331 155147 18379 155175
rect 18069 155113 18379 155147
rect 18069 155085 18117 155113
rect 18145 155085 18179 155113
rect 18207 155085 18241 155113
rect 18269 155085 18303 155113
rect 18331 155085 18379 155113
rect 18069 155051 18379 155085
rect 18069 155023 18117 155051
rect 18145 155023 18179 155051
rect 18207 155023 18241 155051
rect 18269 155023 18303 155051
rect 18331 155023 18379 155051
rect 18069 154989 18379 155023
rect 18069 154961 18117 154989
rect 18145 154961 18179 154989
rect 18207 154961 18241 154989
rect 18269 154961 18303 154989
rect 18331 154961 18379 154989
rect 18069 146175 18379 154961
rect 18069 146147 18117 146175
rect 18145 146147 18179 146175
rect 18207 146147 18241 146175
rect 18269 146147 18303 146175
rect 18331 146147 18379 146175
rect 18069 146113 18379 146147
rect 18069 146085 18117 146113
rect 18145 146085 18179 146113
rect 18207 146085 18241 146113
rect 18269 146085 18303 146113
rect 18331 146085 18379 146113
rect 18069 146051 18379 146085
rect 18069 146023 18117 146051
rect 18145 146023 18179 146051
rect 18207 146023 18241 146051
rect 18269 146023 18303 146051
rect 18331 146023 18379 146051
rect 18069 145989 18379 146023
rect 18069 145961 18117 145989
rect 18145 145961 18179 145989
rect 18207 145961 18241 145989
rect 18269 145961 18303 145989
rect 18331 145961 18379 145989
rect 4569 140147 4617 140175
rect 4645 140147 4679 140175
rect 4707 140147 4741 140175
rect 4769 140147 4803 140175
rect 4831 140147 4879 140175
rect 4569 140113 4879 140147
rect 4569 140085 4617 140113
rect 4645 140085 4679 140113
rect 4707 140085 4741 140113
rect 4769 140085 4803 140113
rect 4831 140085 4879 140113
rect 4569 140051 4879 140085
rect 4569 140023 4617 140051
rect 4645 140023 4679 140051
rect 4707 140023 4741 140051
rect 4769 140023 4803 140051
rect 4831 140023 4879 140051
rect 4569 139989 4879 140023
rect 4569 139961 4617 139989
rect 4645 139961 4679 139989
rect 4707 139961 4741 139989
rect 4769 139961 4803 139989
rect 4831 139961 4879 139989
rect 3990 139874 4018 139879
rect 3934 139314 3962 139319
rect 3878 137634 3906 137639
rect 3822 135394 3850 135399
rect 3150 103161 3178 103166
rect 3766 134274 3794 134279
rect 3094 39657 3122 39662
rect 2709 38147 2757 38175
rect 2785 38147 2819 38175
rect 2847 38147 2881 38175
rect 2909 38147 2943 38175
rect 2971 38147 3019 38175
rect 2709 38113 3019 38147
rect 2709 38085 2757 38113
rect 2785 38085 2819 38113
rect 2847 38085 2881 38113
rect 2909 38085 2943 38113
rect 2971 38085 3019 38113
rect 2709 38051 3019 38085
rect 2709 38023 2757 38051
rect 2785 38023 2819 38051
rect 2847 38023 2881 38051
rect 2909 38023 2943 38051
rect 2971 38023 3019 38051
rect 2709 37989 3019 38023
rect 2709 37961 2757 37989
rect 2785 37961 2819 37989
rect 2847 37961 2881 37989
rect 2909 37961 2943 37989
rect 2971 37961 3019 37989
rect 2709 29175 3019 37961
rect 2709 29147 2757 29175
rect 2785 29147 2819 29175
rect 2847 29147 2881 29175
rect 2909 29147 2943 29175
rect 2971 29147 3019 29175
rect 2709 29113 3019 29147
rect 2709 29085 2757 29113
rect 2785 29085 2819 29113
rect 2847 29085 2881 29113
rect 2909 29085 2943 29113
rect 2971 29085 3019 29113
rect 2709 29051 3019 29085
rect 2709 29023 2757 29051
rect 2785 29023 2819 29051
rect 2847 29023 2881 29051
rect 2909 29023 2943 29051
rect 2971 29023 3019 29051
rect 2709 28989 3019 29023
rect 2709 28961 2757 28989
rect 2785 28961 2819 28989
rect 2847 28961 2881 28989
rect 2909 28961 2943 28989
rect 2971 28961 3019 28989
rect 2709 20175 3019 28961
rect 2709 20147 2757 20175
rect 2785 20147 2819 20175
rect 2847 20147 2881 20175
rect 2909 20147 2943 20175
rect 2971 20147 3019 20175
rect 2709 20113 3019 20147
rect 2709 20085 2757 20113
rect 2785 20085 2819 20113
rect 2847 20085 2881 20113
rect 2909 20085 2943 20113
rect 2971 20085 3019 20113
rect 2709 20051 3019 20085
rect 2709 20023 2757 20051
rect 2785 20023 2819 20051
rect 2847 20023 2881 20051
rect 2909 20023 2943 20051
rect 2971 20023 3019 20051
rect 2709 19989 3019 20023
rect 2709 19961 2757 19989
rect 2785 19961 2819 19989
rect 2847 19961 2881 19989
rect 2909 19961 2943 19989
rect 2971 19961 3019 19989
rect 2086 4377 2114 4382
rect 2709 11175 3019 19961
rect 3766 18466 3794 134246
rect 3822 32634 3850 135366
rect 3878 60858 3906 137606
rect 3934 82026 3962 139286
rect 3990 89026 4018 139846
rect 3990 88993 4018 88998
rect 4569 131175 4879 139961
rect 6286 140434 6314 140439
rect 4569 131147 4617 131175
rect 4645 131147 4679 131175
rect 4707 131147 4741 131175
rect 4769 131147 4803 131175
rect 4831 131147 4879 131175
rect 4569 131113 4879 131147
rect 4569 131085 4617 131113
rect 4645 131085 4679 131113
rect 4707 131085 4741 131113
rect 4769 131085 4803 131113
rect 4831 131085 4879 131113
rect 4569 131051 4879 131085
rect 4569 131023 4617 131051
rect 4645 131023 4679 131051
rect 4707 131023 4741 131051
rect 4769 131023 4803 131051
rect 4831 131023 4879 131051
rect 4569 130989 4879 131023
rect 4569 130961 4617 130989
rect 4645 130961 4679 130989
rect 4707 130961 4741 130989
rect 4769 130961 4803 130989
rect 4831 130961 4879 130989
rect 4569 122175 4879 130961
rect 4569 122147 4617 122175
rect 4645 122147 4679 122175
rect 4707 122147 4741 122175
rect 4769 122147 4803 122175
rect 4831 122147 4879 122175
rect 4569 122113 4879 122147
rect 4569 122085 4617 122113
rect 4645 122085 4679 122113
rect 4707 122085 4741 122113
rect 4769 122085 4803 122113
rect 4831 122085 4879 122113
rect 4569 122051 4879 122085
rect 4569 122023 4617 122051
rect 4645 122023 4679 122051
rect 4707 122023 4741 122051
rect 4769 122023 4803 122051
rect 4831 122023 4879 122051
rect 4569 121989 4879 122023
rect 4569 121961 4617 121989
rect 4645 121961 4679 121989
rect 4707 121961 4741 121989
rect 4769 121961 4803 121989
rect 4831 121961 4879 121989
rect 4569 113175 4879 121961
rect 4569 113147 4617 113175
rect 4645 113147 4679 113175
rect 4707 113147 4741 113175
rect 4769 113147 4803 113175
rect 4831 113147 4879 113175
rect 4569 113113 4879 113147
rect 4569 113085 4617 113113
rect 4645 113085 4679 113113
rect 4707 113085 4741 113113
rect 4769 113085 4803 113113
rect 4831 113085 4879 113113
rect 4569 113051 4879 113085
rect 4569 113023 4617 113051
rect 4645 113023 4679 113051
rect 4707 113023 4741 113051
rect 4769 113023 4803 113051
rect 4831 113023 4879 113051
rect 4569 112989 4879 113023
rect 4569 112961 4617 112989
rect 4645 112961 4679 112989
rect 4707 112961 4741 112989
rect 4769 112961 4803 112989
rect 4831 112961 4879 112989
rect 4569 104175 4879 112961
rect 4569 104147 4617 104175
rect 4645 104147 4679 104175
rect 4707 104147 4741 104175
rect 4769 104147 4803 104175
rect 4831 104147 4879 104175
rect 4569 104113 4879 104147
rect 4569 104085 4617 104113
rect 4645 104085 4679 104113
rect 4707 104085 4741 104113
rect 4769 104085 4803 104113
rect 4831 104085 4879 104113
rect 4569 104051 4879 104085
rect 4569 104023 4617 104051
rect 4645 104023 4679 104051
rect 4707 104023 4741 104051
rect 4769 104023 4803 104051
rect 4831 104023 4879 104051
rect 4569 103989 4879 104023
rect 4569 103961 4617 103989
rect 4645 103961 4679 103989
rect 4707 103961 4741 103989
rect 4769 103961 4803 103989
rect 4831 103961 4879 103989
rect 4569 95175 4879 103961
rect 4569 95147 4617 95175
rect 4645 95147 4679 95175
rect 4707 95147 4741 95175
rect 4769 95147 4803 95175
rect 4831 95147 4879 95175
rect 4569 95113 4879 95147
rect 4569 95085 4617 95113
rect 4645 95085 4679 95113
rect 4707 95085 4741 95113
rect 4769 95085 4803 95113
rect 4831 95085 4879 95113
rect 4569 95051 4879 95085
rect 4569 95023 4617 95051
rect 4645 95023 4679 95051
rect 4707 95023 4741 95051
rect 4769 95023 4803 95051
rect 4831 95023 4879 95051
rect 4569 94989 4879 95023
rect 4569 94961 4617 94989
rect 4645 94961 4679 94989
rect 4707 94961 4741 94989
rect 4769 94961 4803 94989
rect 4831 94961 4879 94989
rect 3934 81993 3962 81998
rect 4569 86175 4879 94961
rect 4569 86147 4617 86175
rect 4645 86147 4679 86175
rect 4707 86147 4741 86175
rect 4769 86147 4803 86175
rect 4831 86147 4879 86175
rect 4569 86113 4879 86147
rect 4569 86085 4617 86113
rect 4645 86085 4679 86113
rect 4707 86085 4741 86113
rect 4769 86085 4803 86113
rect 4831 86085 4879 86113
rect 4569 86051 4879 86085
rect 4569 86023 4617 86051
rect 4645 86023 4679 86051
rect 4707 86023 4741 86051
rect 4769 86023 4803 86051
rect 4831 86023 4879 86051
rect 4569 85989 4879 86023
rect 4569 85961 4617 85989
rect 4645 85961 4679 85989
rect 4707 85961 4741 85989
rect 4769 85961 4803 85989
rect 4831 85961 4879 85989
rect 3878 60825 3906 60830
rect 4569 77175 4879 85961
rect 4569 77147 4617 77175
rect 4645 77147 4679 77175
rect 4707 77147 4741 77175
rect 4769 77147 4803 77175
rect 4831 77147 4879 77175
rect 4569 77113 4879 77147
rect 4569 77085 4617 77113
rect 4645 77085 4679 77113
rect 4707 77085 4741 77113
rect 4769 77085 4803 77113
rect 4831 77085 4879 77113
rect 4569 77051 4879 77085
rect 4569 77023 4617 77051
rect 4645 77023 4679 77051
rect 4707 77023 4741 77051
rect 4769 77023 4803 77051
rect 4831 77023 4879 77051
rect 4569 76989 4879 77023
rect 4569 76961 4617 76989
rect 4645 76961 4679 76989
rect 4707 76961 4741 76989
rect 4769 76961 4803 76989
rect 4831 76961 4879 76989
rect 4569 68175 4879 76961
rect 4569 68147 4617 68175
rect 4645 68147 4679 68175
rect 4707 68147 4741 68175
rect 4769 68147 4803 68175
rect 4831 68147 4879 68175
rect 4569 68113 4879 68147
rect 4569 68085 4617 68113
rect 4645 68085 4679 68113
rect 4707 68085 4741 68113
rect 4769 68085 4803 68113
rect 4831 68085 4879 68113
rect 4569 68051 4879 68085
rect 4569 68023 4617 68051
rect 4645 68023 4679 68051
rect 4707 68023 4741 68051
rect 4769 68023 4803 68051
rect 4831 68023 4879 68051
rect 4569 67989 4879 68023
rect 4569 67961 4617 67989
rect 4645 67961 4679 67989
rect 4707 67961 4741 67989
rect 4769 67961 4803 67989
rect 4831 67961 4879 67989
rect 3822 32601 3850 32606
rect 4569 59175 4879 67961
rect 4569 59147 4617 59175
rect 4645 59147 4679 59175
rect 4707 59147 4741 59175
rect 4769 59147 4803 59175
rect 4831 59147 4879 59175
rect 4569 59113 4879 59147
rect 4569 59085 4617 59113
rect 4645 59085 4679 59113
rect 4707 59085 4741 59113
rect 4769 59085 4803 59113
rect 4831 59085 4879 59113
rect 4569 59051 4879 59085
rect 4569 59023 4617 59051
rect 4645 59023 4679 59051
rect 4707 59023 4741 59051
rect 4769 59023 4803 59051
rect 4831 59023 4879 59051
rect 4569 58989 4879 59023
rect 4569 58961 4617 58989
rect 4645 58961 4679 58989
rect 4707 58961 4741 58989
rect 4769 58961 4803 58989
rect 4831 58961 4879 58989
rect 4569 50175 4879 58961
rect 4569 50147 4617 50175
rect 4645 50147 4679 50175
rect 4707 50147 4741 50175
rect 4769 50147 4803 50175
rect 4831 50147 4879 50175
rect 4569 50113 4879 50147
rect 4569 50085 4617 50113
rect 4645 50085 4679 50113
rect 4707 50085 4741 50113
rect 4769 50085 4803 50113
rect 4831 50085 4879 50113
rect 4569 50051 4879 50085
rect 4569 50023 4617 50051
rect 4645 50023 4679 50051
rect 4707 50023 4741 50051
rect 4769 50023 4803 50051
rect 4831 50023 4879 50051
rect 4569 49989 4879 50023
rect 4569 49961 4617 49989
rect 4645 49961 4679 49989
rect 4707 49961 4741 49989
rect 4769 49961 4803 49989
rect 4831 49961 4879 49989
rect 4569 41175 4879 49961
rect 4569 41147 4617 41175
rect 4645 41147 4679 41175
rect 4707 41147 4741 41175
rect 4769 41147 4803 41175
rect 4831 41147 4879 41175
rect 4569 41113 4879 41147
rect 4569 41085 4617 41113
rect 4645 41085 4679 41113
rect 4707 41085 4741 41113
rect 4769 41085 4803 41113
rect 4831 41085 4879 41113
rect 4569 41051 4879 41085
rect 4569 41023 4617 41051
rect 4645 41023 4679 41051
rect 4707 41023 4741 41051
rect 4769 41023 4803 41051
rect 4831 41023 4879 41051
rect 4569 40989 4879 41023
rect 4569 40961 4617 40989
rect 4645 40961 4679 40989
rect 4707 40961 4741 40989
rect 4769 40961 4803 40989
rect 4831 40961 4879 40989
rect 3766 18433 3794 18438
rect 4569 32175 4879 40961
rect 4569 32147 4617 32175
rect 4645 32147 4679 32175
rect 4707 32147 4741 32175
rect 4769 32147 4803 32175
rect 4831 32147 4879 32175
rect 4569 32113 4879 32147
rect 4569 32085 4617 32113
rect 4645 32085 4679 32113
rect 4707 32085 4741 32113
rect 4769 32085 4803 32113
rect 4831 32085 4879 32113
rect 4569 32051 4879 32085
rect 4569 32023 4617 32051
rect 4645 32023 4679 32051
rect 4707 32023 4741 32051
rect 4769 32023 4803 32051
rect 4831 32023 4879 32051
rect 4569 31989 4879 32023
rect 4569 31961 4617 31989
rect 4645 31961 4679 31989
rect 4707 31961 4741 31989
rect 4769 31961 4803 31989
rect 4831 31961 4879 31989
rect 4569 23175 4879 31961
rect 5446 134834 5474 134839
rect 5446 25578 5474 134806
rect 6286 96026 6314 140406
rect 6286 95993 6314 95998
rect 7126 138754 7154 138759
rect 7126 74858 7154 138726
rect 18069 137175 18379 145961
rect 18069 137147 18117 137175
rect 18145 137147 18179 137175
rect 18207 137147 18241 137175
rect 18269 137147 18303 137175
rect 18331 137147 18379 137175
rect 18069 137113 18379 137147
rect 18069 137085 18117 137113
rect 18145 137085 18179 137113
rect 18207 137085 18241 137113
rect 18269 137085 18303 137113
rect 18331 137085 18379 137113
rect 18069 137051 18379 137085
rect 18069 137023 18117 137051
rect 18145 137023 18179 137051
rect 18207 137023 18241 137051
rect 18269 137023 18303 137051
rect 18331 137023 18379 137051
rect 18069 136989 18379 137023
rect 18069 136961 18117 136989
rect 18145 136961 18179 136989
rect 18207 136961 18241 136989
rect 18269 136961 18303 136989
rect 18331 136961 18379 136989
rect 18069 128175 18379 136961
rect 19929 167175 20239 170745
rect 19929 167147 19977 167175
rect 20005 167147 20039 167175
rect 20067 167147 20101 167175
rect 20129 167147 20163 167175
rect 20191 167147 20239 167175
rect 19929 167113 20239 167147
rect 19929 167085 19977 167113
rect 20005 167085 20039 167113
rect 20067 167085 20101 167113
rect 20129 167085 20163 167113
rect 20191 167085 20239 167113
rect 19929 167051 20239 167085
rect 19929 167023 19977 167051
rect 20005 167023 20039 167051
rect 20067 167023 20101 167051
rect 20129 167023 20163 167051
rect 20191 167023 20239 167051
rect 19929 166989 20239 167023
rect 19929 166961 19977 166989
rect 20005 166961 20039 166989
rect 20067 166961 20101 166989
rect 20129 166961 20163 166989
rect 20191 166961 20239 166989
rect 19929 158175 20239 166961
rect 19929 158147 19977 158175
rect 20005 158147 20039 158175
rect 20067 158147 20101 158175
rect 20129 158147 20163 158175
rect 20191 158147 20239 158175
rect 19929 158113 20239 158147
rect 19929 158085 19977 158113
rect 20005 158085 20039 158113
rect 20067 158085 20101 158113
rect 20129 158085 20163 158113
rect 20191 158085 20239 158113
rect 19929 158051 20239 158085
rect 19929 158023 19977 158051
rect 20005 158023 20039 158051
rect 20067 158023 20101 158051
rect 20129 158023 20163 158051
rect 20191 158023 20239 158051
rect 19929 157989 20239 158023
rect 19929 157961 19977 157989
rect 20005 157961 20039 157989
rect 20067 157961 20101 157989
rect 20129 157961 20163 157989
rect 20191 157961 20239 157989
rect 19929 149175 20239 157961
rect 33429 164175 33739 170745
rect 33429 164147 33477 164175
rect 33505 164147 33539 164175
rect 33567 164147 33601 164175
rect 33629 164147 33663 164175
rect 33691 164147 33739 164175
rect 33429 164113 33739 164147
rect 33429 164085 33477 164113
rect 33505 164085 33539 164113
rect 33567 164085 33601 164113
rect 33629 164085 33663 164113
rect 33691 164085 33739 164113
rect 33429 164051 33739 164085
rect 33429 164023 33477 164051
rect 33505 164023 33539 164051
rect 33567 164023 33601 164051
rect 33629 164023 33663 164051
rect 33691 164023 33739 164051
rect 33429 163989 33739 164023
rect 33429 163961 33477 163989
rect 33505 163961 33539 163989
rect 33567 163961 33601 163989
rect 33629 163961 33663 163989
rect 33691 163961 33739 163989
rect 32224 155175 32384 155192
rect 32224 155147 32259 155175
rect 32287 155147 32321 155175
rect 32349 155147 32384 155175
rect 32224 155113 32384 155147
rect 32224 155085 32259 155113
rect 32287 155085 32321 155113
rect 32349 155085 32384 155113
rect 32224 155051 32384 155085
rect 32224 155023 32259 155051
rect 32287 155023 32321 155051
rect 32349 155023 32384 155051
rect 32224 154989 32384 155023
rect 32224 154961 32259 154989
rect 32287 154961 32321 154989
rect 32349 154961 32384 154989
rect 32224 154944 32384 154961
rect 33429 155175 33739 163961
rect 33429 155147 33477 155175
rect 33505 155147 33539 155175
rect 33567 155147 33601 155175
rect 33629 155147 33663 155175
rect 33691 155147 33739 155175
rect 33429 155113 33739 155147
rect 33429 155085 33477 155113
rect 33505 155085 33539 155113
rect 33567 155085 33601 155113
rect 33629 155085 33663 155113
rect 33691 155085 33739 155113
rect 33429 155051 33739 155085
rect 33429 155023 33477 155051
rect 33505 155023 33539 155051
rect 33567 155023 33601 155051
rect 33629 155023 33663 155051
rect 33691 155023 33739 155051
rect 33429 154989 33739 155023
rect 33429 154961 33477 154989
rect 33505 154961 33539 154989
rect 33567 154961 33601 154989
rect 33629 154961 33663 154989
rect 33691 154961 33739 154989
rect 19929 149147 19977 149175
rect 20005 149147 20039 149175
rect 20067 149147 20101 149175
rect 20129 149147 20163 149175
rect 20191 149147 20239 149175
rect 19929 149113 20239 149147
rect 19929 149085 19977 149113
rect 20005 149085 20039 149113
rect 20067 149085 20101 149113
rect 20129 149085 20163 149113
rect 20191 149085 20239 149113
rect 19929 149051 20239 149085
rect 19929 149023 19977 149051
rect 20005 149023 20039 149051
rect 20067 149023 20101 149051
rect 20129 149023 20163 149051
rect 20191 149023 20239 149051
rect 19929 148989 20239 149023
rect 19929 148961 19977 148989
rect 20005 148961 20039 148989
rect 20067 148961 20101 148989
rect 20129 148961 20163 148989
rect 20191 148961 20239 148989
rect 19929 140175 20239 148961
rect 32224 146175 32384 146192
rect 32224 146147 32259 146175
rect 32287 146147 32321 146175
rect 32349 146147 32384 146175
rect 32224 146113 32384 146147
rect 32224 146085 32259 146113
rect 32287 146085 32321 146113
rect 32349 146085 32384 146113
rect 32224 146051 32384 146085
rect 32224 146023 32259 146051
rect 32287 146023 32321 146051
rect 32349 146023 32384 146051
rect 32224 145989 32384 146023
rect 32224 145961 32259 145989
rect 32287 145961 32321 145989
rect 32349 145961 32384 145989
rect 32224 145944 32384 145961
rect 33429 146175 33739 154961
rect 33429 146147 33477 146175
rect 33505 146147 33539 146175
rect 33567 146147 33601 146175
rect 33629 146147 33663 146175
rect 33691 146147 33739 146175
rect 33429 146113 33739 146147
rect 33429 146085 33477 146113
rect 33505 146085 33539 146113
rect 33567 146085 33601 146113
rect 33629 146085 33663 146113
rect 33691 146085 33739 146113
rect 33429 146051 33739 146085
rect 33429 146023 33477 146051
rect 33505 146023 33539 146051
rect 33567 146023 33601 146051
rect 33629 146023 33663 146051
rect 33691 146023 33739 146051
rect 33429 145989 33739 146023
rect 33429 145961 33477 145989
rect 33505 145961 33539 145989
rect 33567 145961 33601 145989
rect 33629 145961 33663 145989
rect 33691 145961 33739 145989
rect 28238 143234 28266 143239
rect 28182 142674 28210 142679
rect 19929 140147 19977 140175
rect 20005 140147 20039 140175
rect 20067 140147 20101 140175
rect 20129 140147 20163 140175
rect 20191 140147 20239 140175
rect 19929 140113 20239 140147
rect 19929 140085 19977 140113
rect 20005 140085 20039 140113
rect 20067 140085 20101 140113
rect 20129 140085 20163 140113
rect 20191 140085 20239 140113
rect 19929 140051 20239 140085
rect 19929 140023 19977 140051
rect 20005 140023 20039 140051
rect 20067 140023 20101 140051
rect 20129 140023 20163 140051
rect 20191 140023 20239 140051
rect 19929 139989 20239 140023
rect 19929 139961 19977 139989
rect 20005 139961 20039 139989
rect 20067 139961 20101 139989
rect 20129 139961 20163 139989
rect 20191 139961 20239 139989
rect 18069 128147 18117 128175
rect 18145 128147 18179 128175
rect 18207 128147 18241 128175
rect 18269 128147 18303 128175
rect 18331 128147 18379 128175
rect 18069 128113 18379 128147
rect 18069 128085 18117 128113
rect 18145 128085 18179 128113
rect 18207 128085 18241 128113
rect 18269 128085 18303 128113
rect 18331 128085 18379 128113
rect 18069 128051 18379 128085
rect 18069 128023 18117 128051
rect 18145 128023 18179 128051
rect 18207 128023 18241 128051
rect 18269 128023 18303 128051
rect 18331 128023 18379 128051
rect 18069 127989 18379 128023
rect 18069 127961 18117 127989
rect 18145 127961 18179 127989
rect 18207 127961 18241 127989
rect 18269 127961 18303 127989
rect 18331 127961 18379 127989
rect 18069 119175 18379 127961
rect 18069 119147 18117 119175
rect 18145 119147 18179 119175
rect 18207 119147 18241 119175
rect 18269 119147 18303 119175
rect 18331 119147 18379 119175
rect 18069 119113 18379 119147
rect 18069 119085 18117 119113
rect 18145 119085 18179 119113
rect 18207 119085 18241 119113
rect 18269 119085 18303 119113
rect 18331 119085 18379 119113
rect 18069 119051 18379 119085
rect 18069 119023 18117 119051
rect 18145 119023 18179 119051
rect 18207 119023 18241 119051
rect 18269 119023 18303 119051
rect 18331 119023 18379 119051
rect 18069 118989 18379 119023
rect 18069 118961 18117 118989
rect 18145 118961 18179 118989
rect 18207 118961 18241 118989
rect 18269 118961 18303 118989
rect 18331 118961 18379 118989
rect 18069 110175 18379 118961
rect 18069 110147 18117 110175
rect 18145 110147 18179 110175
rect 18207 110147 18241 110175
rect 18269 110147 18303 110175
rect 18331 110147 18379 110175
rect 18069 110113 18379 110147
rect 18069 110085 18117 110113
rect 18145 110085 18179 110113
rect 18207 110085 18241 110113
rect 18269 110085 18303 110113
rect 18331 110085 18379 110113
rect 18069 110051 18379 110085
rect 18069 110023 18117 110051
rect 18145 110023 18179 110051
rect 18207 110023 18241 110051
rect 18269 110023 18303 110051
rect 18331 110023 18379 110051
rect 18069 109989 18379 110023
rect 18069 109961 18117 109989
rect 18145 109961 18179 109989
rect 18207 109961 18241 109989
rect 18269 109961 18303 109989
rect 18331 109961 18379 109989
rect 16224 101175 16384 101192
rect 16224 101147 16259 101175
rect 16287 101147 16321 101175
rect 16349 101147 16384 101175
rect 16224 101113 16384 101147
rect 16224 101085 16259 101113
rect 16287 101085 16321 101113
rect 16349 101085 16384 101113
rect 16224 101051 16384 101085
rect 16224 101023 16259 101051
rect 16287 101023 16321 101051
rect 16349 101023 16384 101051
rect 16224 100989 16384 101023
rect 16224 100961 16259 100989
rect 16287 100961 16321 100989
rect 16349 100961 16384 100989
rect 16224 100944 16384 100961
rect 18069 101175 18379 109961
rect 18069 101147 18117 101175
rect 18145 101147 18179 101175
rect 18207 101147 18241 101175
rect 18269 101147 18303 101175
rect 18331 101147 18379 101175
rect 18069 101113 18379 101147
rect 18069 101085 18117 101113
rect 18145 101085 18179 101113
rect 18207 101085 18241 101113
rect 18269 101085 18303 101113
rect 18331 101085 18379 101113
rect 18069 101051 18379 101085
rect 18069 101023 18117 101051
rect 18145 101023 18179 101051
rect 18207 101023 18241 101051
rect 18269 101023 18303 101051
rect 18331 101023 18379 101051
rect 18069 100989 18379 101023
rect 18069 100961 18117 100989
rect 18145 100961 18179 100989
rect 18207 100961 18241 100989
rect 18269 100961 18303 100989
rect 18331 100961 18379 100989
rect 16224 92175 16384 92192
rect 16224 92147 16259 92175
rect 16287 92147 16321 92175
rect 16349 92147 16384 92175
rect 16224 92113 16384 92147
rect 16224 92085 16259 92113
rect 16287 92085 16321 92113
rect 16349 92085 16384 92113
rect 16224 92051 16384 92085
rect 16224 92023 16259 92051
rect 16287 92023 16321 92051
rect 16349 92023 16384 92051
rect 16224 91989 16384 92023
rect 16224 91961 16259 91989
rect 16287 91961 16321 91989
rect 16349 91961 16384 91989
rect 16224 91944 16384 91961
rect 18069 92175 18379 100961
rect 18069 92147 18117 92175
rect 18145 92147 18179 92175
rect 18207 92147 18241 92175
rect 18269 92147 18303 92175
rect 18331 92147 18379 92175
rect 18069 92113 18379 92147
rect 18069 92085 18117 92113
rect 18145 92085 18179 92113
rect 18207 92085 18241 92113
rect 18269 92085 18303 92113
rect 18331 92085 18379 92113
rect 18069 92051 18379 92085
rect 18069 92023 18117 92051
rect 18145 92023 18179 92051
rect 18207 92023 18241 92051
rect 18269 92023 18303 92051
rect 18331 92023 18379 92051
rect 18069 91989 18379 92023
rect 18069 91961 18117 91989
rect 18145 91961 18179 91989
rect 18207 91961 18241 91989
rect 18269 91961 18303 91989
rect 18331 91961 18379 91989
rect 16224 83175 16384 83192
rect 16224 83147 16259 83175
rect 16287 83147 16321 83175
rect 16349 83147 16384 83175
rect 16224 83113 16384 83147
rect 16224 83085 16259 83113
rect 16287 83085 16321 83113
rect 16349 83085 16384 83113
rect 16224 83051 16384 83085
rect 16224 83023 16259 83051
rect 16287 83023 16321 83051
rect 16349 83023 16384 83051
rect 16224 82989 16384 83023
rect 16224 82961 16259 82989
rect 16287 82961 16321 82989
rect 16349 82961 16384 82989
rect 16224 82944 16384 82961
rect 18069 83175 18379 91961
rect 18069 83147 18117 83175
rect 18145 83147 18179 83175
rect 18207 83147 18241 83175
rect 18269 83147 18303 83175
rect 18331 83147 18379 83175
rect 18069 83113 18379 83147
rect 18069 83085 18117 83113
rect 18145 83085 18179 83113
rect 18207 83085 18241 83113
rect 18269 83085 18303 83113
rect 18331 83085 18379 83113
rect 18069 83051 18379 83085
rect 18069 83023 18117 83051
rect 18145 83023 18179 83051
rect 18207 83023 18241 83051
rect 18269 83023 18303 83051
rect 18331 83023 18379 83051
rect 18069 82989 18379 83023
rect 18069 82961 18117 82989
rect 18145 82961 18179 82989
rect 18207 82961 18241 82989
rect 18269 82961 18303 82989
rect 18331 82961 18379 82989
rect 7126 74825 7154 74830
rect 5446 25545 5474 25550
rect 18069 74175 18379 82961
rect 19278 132034 19306 132039
rect 19278 75362 19306 132006
rect 19278 75138 19306 75334
rect 19278 75105 19306 75110
rect 19929 131175 20239 139961
rect 28126 141554 28154 141559
rect 19929 131147 19977 131175
rect 20005 131147 20039 131175
rect 20067 131147 20101 131175
rect 20129 131147 20163 131175
rect 20191 131147 20239 131175
rect 19929 131113 20239 131147
rect 19929 131085 19977 131113
rect 20005 131085 20039 131113
rect 20067 131085 20101 131113
rect 20129 131085 20163 131113
rect 20191 131085 20239 131113
rect 19929 131051 20239 131085
rect 19929 131023 19977 131051
rect 20005 131023 20039 131051
rect 20067 131023 20101 131051
rect 20129 131023 20163 131051
rect 20191 131023 20239 131051
rect 19929 130989 20239 131023
rect 19929 130961 19977 130989
rect 20005 130961 20039 130989
rect 20067 130961 20101 130989
rect 20129 130961 20163 130989
rect 20191 130961 20239 130989
rect 19929 122175 20239 130961
rect 19929 122147 19977 122175
rect 20005 122147 20039 122175
rect 20067 122147 20101 122175
rect 20129 122147 20163 122175
rect 20191 122147 20239 122175
rect 19929 122113 20239 122147
rect 19929 122085 19977 122113
rect 20005 122085 20039 122113
rect 20067 122085 20101 122113
rect 20129 122085 20163 122113
rect 20191 122085 20239 122113
rect 19929 122051 20239 122085
rect 19929 122023 19977 122051
rect 20005 122023 20039 122051
rect 20067 122023 20101 122051
rect 20129 122023 20163 122051
rect 20191 122023 20239 122051
rect 19929 121989 20239 122023
rect 19929 121961 19977 121989
rect 20005 121961 20039 121989
rect 20067 121961 20101 121989
rect 20129 121961 20163 121989
rect 20191 121961 20239 121989
rect 19929 113175 20239 121961
rect 19929 113147 19977 113175
rect 20005 113147 20039 113175
rect 20067 113147 20101 113175
rect 20129 113147 20163 113175
rect 20191 113147 20239 113175
rect 19929 113113 20239 113147
rect 19929 113085 19977 113113
rect 20005 113085 20039 113113
rect 20067 113085 20101 113113
rect 20129 113085 20163 113113
rect 20191 113085 20239 113113
rect 19929 113051 20239 113085
rect 19929 113023 19977 113051
rect 20005 113023 20039 113051
rect 20067 113023 20101 113051
rect 20129 113023 20163 113051
rect 20191 113023 20239 113051
rect 19929 112989 20239 113023
rect 19929 112961 19977 112989
rect 20005 112961 20039 112989
rect 20067 112961 20101 112989
rect 20129 112961 20163 112989
rect 20191 112961 20239 112989
rect 19929 104175 20239 112961
rect 19929 104147 19977 104175
rect 20005 104147 20039 104175
rect 20067 104147 20101 104175
rect 20129 104147 20163 104175
rect 20191 104147 20239 104175
rect 19929 104113 20239 104147
rect 19929 104085 19977 104113
rect 20005 104085 20039 104113
rect 20067 104085 20101 104113
rect 20129 104085 20163 104113
rect 20191 104085 20239 104113
rect 19929 104051 20239 104085
rect 19929 104023 19977 104051
rect 20005 104023 20039 104051
rect 20067 104023 20101 104051
rect 20129 104023 20163 104051
rect 20191 104023 20239 104051
rect 19929 103989 20239 104023
rect 19929 103961 19977 103989
rect 20005 103961 20039 103989
rect 20067 103961 20101 103989
rect 20129 103961 20163 103989
rect 20191 103961 20239 103989
rect 19929 95175 20239 103961
rect 19929 95147 19977 95175
rect 20005 95147 20039 95175
rect 20067 95147 20101 95175
rect 20129 95147 20163 95175
rect 20191 95147 20239 95175
rect 19929 95113 20239 95147
rect 19929 95085 19977 95113
rect 20005 95085 20039 95113
rect 20067 95085 20101 95113
rect 20129 95085 20163 95113
rect 20191 95085 20239 95113
rect 19929 95051 20239 95085
rect 19929 95023 19977 95051
rect 20005 95023 20039 95051
rect 20067 95023 20101 95051
rect 20129 95023 20163 95051
rect 20191 95023 20239 95051
rect 19929 94989 20239 95023
rect 19929 94961 19977 94989
rect 20005 94961 20039 94989
rect 20067 94961 20101 94989
rect 20129 94961 20163 94989
rect 20191 94961 20239 94989
rect 19929 86175 20239 94961
rect 19929 86147 19977 86175
rect 20005 86147 20039 86175
rect 20067 86147 20101 86175
rect 20129 86147 20163 86175
rect 20191 86147 20239 86175
rect 19929 86113 20239 86147
rect 19929 86085 19977 86113
rect 20005 86085 20039 86113
rect 20067 86085 20101 86113
rect 20129 86085 20163 86113
rect 20191 86085 20239 86113
rect 19929 86051 20239 86085
rect 19929 86023 19977 86051
rect 20005 86023 20039 86051
rect 20067 86023 20101 86051
rect 20129 86023 20163 86051
rect 20191 86023 20239 86051
rect 19929 85989 20239 86023
rect 19929 85961 19977 85989
rect 20005 85961 20039 85989
rect 20067 85961 20101 85989
rect 20129 85961 20163 85989
rect 20191 85961 20239 85989
rect 19929 77175 20239 85961
rect 19929 77147 19977 77175
rect 20005 77147 20039 77175
rect 20067 77147 20101 77175
rect 20129 77147 20163 77175
rect 20191 77147 20239 77175
rect 19929 77113 20239 77147
rect 19929 77085 19977 77113
rect 20005 77085 20039 77113
rect 20067 77085 20101 77113
rect 20129 77085 20163 77113
rect 20191 77085 20239 77113
rect 19929 77051 20239 77085
rect 19929 77023 19977 77051
rect 20005 77023 20039 77051
rect 20067 77023 20101 77051
rect 20129 77023 20163 77051
rect 20191 77023 20239 77051
rect 19929 76989 20239 77023
rect 19929 76961 19977 76989
rect 20005 76961 20039 76989
rect 20067 76961 20101 76989
rect 20129 76961 20163 76989
rect 20191 76961 20239 76989
rect 18069 74147 18117 74175
rect 18145 74147 18179 74175
rect 18207 74147 18241 74175
rect 18269 74147 18303 74175
rect 18331 74147 18379 74175
rect 18069 74113 18379 74147
rect 18069 74085 18117 74113
rect 18145 74085 18179 74113
rect 18207 74085 18241 74113
rect 18269 74085 18303 74113
rect 18331 74085 18379 74113
rect 18069 74051 18379 74085
rect 18069 74023 18117 74051
rect 18145 74023 18179 74051
rect 18207 74023 18241 74051
rect 18269 74023 18303 74051
rect 18331 74023 18379 74051
rect 18069 73989 18379 74023
rect 18069 73961 18117 73989
rect 18145 73961 18179 73989
rect 18207 73961 18241 73989
rect 18269 73961 18303 73989
rect 18331 73961 18379 73989
rect 18069 65175 18379 73961
rect 18069 65147 18117 65175
rect 18145 65147 18179 65175
rect 18207 65147 18241 65175
rect 18269 65147 18303 65175
rect 18331 65147 18379 65175
rect 18069 65113 18379 65147
rect 18069 65085 18117 65113
rect 18145 65085 18179 65113
rect 18207 65085 18241 65113
rect 18269 65085 18303 65113
rect 18331 65085 18379 65113
rect 18069 65051 18379 65085
rect 18069 65023 18117 65051
rect 18145 65023 18179 65051
rect 18207 65023 18241 65051
rect 18269 65023 18303 65051
rect 18331 65023 18379 65051
rect 18069 64989 18379 65023
rect 18069 64961 18117 64989
rect 18145 64961 18179 64989
rect 18207 64961 18241 64989
rect 18269 64961 18303 64989
rect 18331 64961 18379 64989
rect 18069 56175 18379 64961
rect 18069 56147 18117 56175
rect 18145 56147 18179 56175
rect 18207 56147 18241 56175
rect 18269 56147 18303 56175
rect 18331 56147 18379 56175
rect 18069 56113 18379 56147
rect 18069 56085 18117 56113
rect 18145 56085 18179 56113
rect 18207 56085 18241 56113
rect 18269 56085 18303 56113
rect 18331 56085 18379 56113
rect 18069 56051 18379 56085
rect 18069 56023 18117 56051
rect 18145 56023 18179 56051
rect 18207 56023 18241 56051
rect 18269 56023 18303 56051
rect 18331 56023 18379 56051
rect 18069 55989 18379 56023
rect 18069 55961 18117 55989
rect 18145 55961 18179 55989
rect 18207 55961 18241 55989
rect 18269 55961 18303 55989
rect 18331 55961 18379 55989
rect 18069 47175 18379 55961
rect 18069 47147 18117 47175
rect 18145 47147 18179 47175
rect 18207 47147 18241 47175
rect 18269 47147 18303 47175
rect 18331 47147 18379 47175
rect 18069 47113 18379 47147
rect 18069 47085 18117 47113
rect 18145 47085 18179 47113
rect 18207 47085 18241 47113
rect 18269 47085 18303 47113
rect 18331 47085 18379 47113
rect 18069 47051 18379 47085
rect 18069 47023 18117 47051
rect 18145 47023 18179 47051
rect 18207 47023 18241 47051
rect 18269 47023 18303 47051
rect 18331 47023 18379 47051
rect 18069 46989 18379 47023
rect 18069 46961 18117 46989
rect 18145 46961 18179 46989
rect 18207 46961 18241 46989
rect 18269 46961 18303 46989
rect 18331 46961 18379 46989
rect 18069 38175 18379 46961
rect 18069 38147 18117 38175
rect 18145 38147 18179 38175
rect 18207 38147 18241 38175
rect 18269 38147 18303 38175
rect 18331 38147 18379 38175
rect 18069 38113 18379 38147
rect 18069 38085 18117 38113
rect 18145 38085 18179 38113
rect 18207 38085 18241 38113
rect 18269 38085 18303 38113
rect 18331 38085 18379 38113
rect 18069 38051 18379 38085
rect 18069 38023 18117 38051
rect 18145 38023 18179 38051
rect 18207 38023 18241 38051
rect 18269 38023 18303 38051
rect 18331 38023 18379 38051
rect 18069 37989 18379 38023
rect 18069 37961 18117 37989
rect 18145 37961 18179 37989
rect 18207 37961 18241 37989
rect 18269 37961 18303 37989
rect 18331 37961 18379 37989
rect 18069 29175 18379 37961
rect 18069 29147 18117 29175
rect 18145 29147 18179 29175
rect 18207 29147 18241 29175
rect 18269 29147 18303 29175
rect 18331 29147 18379 29175
rect 18069 29113 18379 29147
rect 18069 29085 18117 29113
rect 18145 29085 18179 29113
rect 18207 29085 18241 29113
rect 18269 29085 18303 29113
rect 18331 29085 18379 29113
rect 18069 29051 18379 29085
rect 18069 29023 18117 29051
rect 18145 29023 18179 29051
rect 18207 29023 18241 29051
rect 18269 29023 18303 29051
rect 18331 29023 18379 29051
rect 18069 28989 18379 29023
rect 18069 28961 18117 28989
rect 18145 28961 18179 28989
rect 18207 28961 18241 28989
rect 18269 28961 18303 28989
rect 18331 28961 18379 28989
rect 4569 23147 4617 23175
rect 4645 23147 4679 23175
rect 4707 23147 4741 23175
rect 4769 23147 4803 23175
rect 4831 23147 4879 23175
rect 4569 23113 4879 23147
rect 4569 23085 4617 23113
rect 4645 23085 4679 23113
rect 4707 23085 4741 23113
rect 4769 23085 4803 23113
rect 4831 23085 4879 23113
rect 4569 23051 4879 23085
rect 4569 23023 4617 23051
rect 4645 23023 4679 23051
rect 4707 23023 4741 23051
rect 4769 23023 4803 23051
rect 4831 23023 4879 23051
rect 4569 22989 4879 23023
rect 4569 22961 4617 22989
rect 4645 22961 4679 22989
rect 4707 22961 4741 22989
rect 4769 22961 4803 22989
rect 4831 22961 4879 22989
rect 2709 11147 2757 11175
rect 2785 11147 2819 11175
rect 2847 11147 2881 11175
rect 2909 11147 2943 11175
rect 2971 11147 3019 11175
rect 2709 11113 3019 11147
rect 2709 11085 2757 11113
rect 2785 11085 2819 11113
rect 2847 11085 2881 11113
rect 2909 11085 2943 11113
rect 2971 11085 3019 11113
rect 2709 11051 3019 11085
rect 2709 11023 2757 11051
rect 2785 11023 2819 11051
rect 2847 11023 2881 11051
rect 2909 11023 2943 11051
rect 2971 11023 3019 11051
rect 2709 10989 3019 11023
rect 2709 10961 2757 10989
rect 2785 10961 2819 10989
rect 2847 10961 2881 10989
rect 2909 10961 2943 10989
rect 2971 10961 3019 10989
rect -478 2147 -430 2175
rect -402 2147 -368 2175
rect -340 2147 -306 2175
rect -278 2147 -244 2175
rect -216 2147 -168 2175
rect -478 2113 -168 2147
rect -478 2085 -430 2113
rect -402 2085 -368 2113
rect -340 2085 -306 2113
rect -278 2085 -244 2113
rect -216 2085 -168 2113
rect -478 2051 -168 2085
rect -478 2023 -430 2051
rect -402 2023 -368 2051
rect -340 2023 -306 2051
rect -278 2023 -244 2051
rect -216 2023 -168 2051
rect -478 1989 -168 2023
rect -478 1961 -430 1989
rect -402 1961 -368 1989
rect -340 1961 -306 1989
rect -278 1961 -244 1989
rect -216 1961 -168 1989
rect -478 -80 -168 1961
rect -478 -108 -430 -80
rect -402 -108 -368 -80
rect -340 -108 -306 -80
rect -278 -108 -244 -80
rect -216 -108 -168 -80
rect -478 -142 -168 -108
rect -478 -170 -430 -142
rect -402 -170 -368 -142
rect -340 -170 -306 -142
rect -278 -170 -244 -142
rect -216 -170 -168 -142
rect -478 -204 -168 -170
rect -478 -232 -430 -204
rect -402 -232 -368 -204
rect -340 -232 -306 -204
rect -278 -232 -244 -204
rect -216 -232 -168 -204
rect -478 -266 -168 -232
rect -478 -294 -430 -266
rect -402 -294 -368 -266
rect -340 -294 -306 -266
rect -278 -294 -244 -266
rect -216 -294 -168 -266
rect -478 -342 -168 -294
rect 2709 2175 3019 10961
rect 2709 2147 2757 2175
rect 2785 2147 2819 2175
rect 2847 2147 2881 2175
rect 2909 2147 2943 2175
rect 2971 2147 3019 2175
rect 2709 2113 3019 2147
rect 2709 2085 2757 2113
rect 2785 2085 2819 2113
rect 2847 2085 2881 2113
rect 2909 2085 2943 2113
rect 2971 2085 3019 2113
rect 2709 2051 3019 2085
rect 2709 2023 2757 2051
rect 2785 2023 2819 2051
rect 2847 2023 2881 2051
rect 2909 2023 2943 2051
rect 2971 2023 3019 2051
rect 2709 1989 3019 2023
rect 2709 1961 2757 1989
rect 2785 1961 2819 1989
rect 2847 1961 2881 1989
rect 2909 1961 2943 1989
rect 2971 1961 3019 1989
rect 2709 -80 3019 1961
rect 2709 -108 2757 -80
rect 2785 -108 2819 -80
rect 2847 -108 2881 -80
rect 2909 -108 2943 -80
rect 2971 -108 3019 -80
rect 2709 -142 3019 -108
rect 2709 -170 2757 -142
rect 2785 -170 2819 -142
rect 2847 -170 2881 -142
rect 2909 -170 2943 -142
rect 2971 -170 3019 -142
rect 2709 -204 3019 -170
rect 2709 -232 2757 -204
rect 2785 -232 2819 -204
rect 2847 -232 2881 -204
rect 2909 -232 2943 -204
rect 2971 -232 3019 -204
rect 2709 -266 3019 -232
rect 2709 -294 2757 -266
rect 2785 -294 2819 -266
rect 2847 -294 2881 -266
rect 2909 -294 2943 -266
rect 2971 -294 3019 -266
rect -958 -588 -910 -560
rect -882 -588 -848 -560
rect -820 -588 -786 -560
rect -758 -588 -724 -560
rect -696 -588 -648 -560
rect -958 -622 -648 -588
rect -958 -650 -910 -622
rect -882 -650 -848 -622
rect -820 -650 -786 -622
rect -758 -650 -724 -622
rect -696 -650 -648 -622
rect -958 -684 -648 -650
rect -958 -712 -910 -684
rect -882 -712 -848 -684
rect -820 -712 -786 -684
rect -758 -712 -724 -684
rect -696 -712 -648 -684
rect -958 -746 -648 -712
rect -958 -774 -910 -746
rect -882 -774 -848 -746
rect -820 -774 -786 -746
rect -758 -774 -724 -746
rect -696 -774 -648 -746
rect -958 -822 -648 -774
rect 2709 -822 3019 -294
rect 4569 14175 4879 22961
rect 4569 14147 4617 14175
rect 4645 14147 4679 14175
rect 4707 14147 4741 14175
rect 4769 14147 4803 14175
rect 4831 14147 4879 14175
rect 4569 14113 4879 14147
rect 4569 14085 4617 14113
rect 4645 14085 4679 14113
rect 4707 14085 4741 14113
rect 4769 14085 4803 14113
rect 4831 14085 4879 14113
rect 4569 14051 4879 14085
rect 4569 14023 4617 14051
rect 4645 14023 4679 14051
rect 4707 14023 4741 14051
rect 4769 14023 4803 14051
rect 4831 14023 4879 14051
rect 4569 13989 4879 14023
rect 4569 13961 4617 13989
rect 4645 13961 4679 13989
rect 4707 13961 4741 13989
rect 4769 13961 4803 13989
rect 4831 13961 4879 13989
rect 4569 5175 4879 13961
rect 4569 5147 4617 5175
rect 4645 5147 4679 5175
rect 4707 5147 4741 5175
rect 4769 5147 4803 5175
rect 4831 5147 4879 5175
rect 4569 5113 4879 5147
rect 4569 5085 4617 5113
rect 4645 5085 4679 5113
rect 4707 5085 4741 5113
rect 4769 5085 4803 5113
rect 4831 5085 4879 5113
rect 4569 5051 4879 5085
rect 4569 5023 4617 5051
rect 4645 5023 4679 5051
rect 4707 5023 4741 5051
rect 4769 5023 4803 5051
rect 4831 5023 4879 5051
rect 4569 4989 4879 5023
rect 4569 4961 4617 4989
rect 4645 4961 4679 4989
rect 4707 4961 4741 4989
rect 4769 4961 4803 4989
rect 4831 4961 4879 4989
rect 4569 -560 4879 4961
rect 4569 -588 4617 -560
rect 4645 -588 4679 -560
rect 4707 -588 4741 -560
rect 4769 -588 4803 -560
rect 4831 -588 4879 -560
rect 4569 -622 4879 -588
rect 4569 -650 4617 -622
rect 4645 -650 4679 -622
rect 4707 -650 4741 -622
rect 4769 -650 4803 -622
rect 4831 -650 4879 -622
rect 4569 -684 4879 -650
rect 4569 -712 4617 -684
rect 4645 -712 4679 -684
rect 4707 -712 4741 -684
rect 4769 -712 4803 -684
rect 4831 -712 4879 -684
rect 4569 -746 4879 -712
rect 4569 -774 4617 -746
rect 4645 -774 4679 -746
rect 4707 -774 4741 -746
rect 4769 -774 4803 -746
rect 4831 -774 4879 -746
rect 4569 -822 4879 -774
rect 18069 20175 18379 28961
rect 18069 20147 18117 20175
rect 18145 20147 18179 20175
rect 18207 20147 18241 20175
rect 18269 20147 18303 20175
rect 18331 20147 18379 20175
rect 18069 20113 18379 20147
rect 18069 20085 18117 20113
rect 18145 20085 18179 20113
rect 18207 20085 18241 20113
rect 18269 20085 18303 20113
rect 18331 20085 18379 20113
rect 18069 20051 18379 20085
rect 18069 20023 18117 20051
rect 18145 20023 18179 20051
rect 18207 20023 18241 20051
rect 18269 20023 18303 20051
rect 18331 20023 18379 20051
rect 18069 19989 18379 20023
rect 18069 19961 18117 19989
rect 18145 19961 18179 19989
rect 18207 19961 18241 19989
rect 18269 19961 18303 19989
rect 18331 19961 18379 19989
rect 18069 11175 18379 19961
rect 18069 11147 18117 11175
rect 18145 11147 18179 11175
rect 18207 11147 18241 11175
rect 18269 11147 18303 11175
rect 18331 11147 18379 11175
rect 18069 11113 18379 11147
rect 18069 11085 18117 11113
rect 18145 11085 18179 11113
rect 18207 11085 18241 11113
rect 18269 11085 18303 11113
rect 18331 11085 18379 11113
rect 18069 11051 18379 11085
rect 18069 11023 18117 11051
rect 18145 11023 18179 11051
rect 18207 11023 18241 11051
rect 18269 11023 18303 11051
rect 18331 11023 18379 11051
rect 18069 10989 18379 11023
rect 18069 10961 18117 10989
rect 18145 10961 18179 10989
rect 18207 10961 18241 10989
rect 18269 10961 18303 10989
rect 18331 10961 18379 10989
rect 18069 2175 18379 10961
rect 18069 2147 18117 2175
rect 18145 2147 18179 2175
rect 18207 2147 18241 2175
rect 18269 2147 18303 2175
rect 18331 2147 18379 2175
rect 18069 2113 18379 2147
rect 18069 2085 18117 2113
rect 18145 2085 18179 2113
rect 18207 2085 18241 2113
rect 18269 2085 18303 2113
rect 18331 2085 18379 2113
rect 18069 2051 18379 2085
rect 18069 2023 18117 2051
rect 18145 2023 18179 2051
rect 18207 2023 18241 2051
rect 18269 2023 18303 2051
rect 18331 2023 18379 2051
rect 18069 1989 18379 2023
rect 18069 1961 18117 1989
rect 18145 1961 18179 1989
rect 18207 1961 18241 1989
rect 18269 1961 18303 1989
rect 18331 1961 18379 1989
rect 18069 -80 18379 1961
rect 18069 -108 18117 -80
rect 18145 -108 18179 -80
rect 18207 -108 18241 -80
rect 18269 -108 18303 -80
rect 18331 -108 18379 -80
rect 18069 -142 18379 -108
rect 18069 -170 18117 -142
rect 18145 -170 18179 -142
rect 18207 -170 18241 -142
rect 18269 -170 18303 -142
rect 18331 -170 18379 -142
rect 18069 -204 18379 -170
rect 18069 -232 18117 -204
rect 18145 -232 18179 -204
rect 18207 -232 18241 -204
rect 18269 -232 18303 -204
rect 18331 -232 18379 -204
rect 18069 -266 18379 -232
rect 18069 -294 18117 -266
rect 18145 -294 18179 -266
rect 18207 -294 18241 -266
rect 18269 -294 18303 -266
rect 18331 -294 18379 -266
rect 18069 -822 18379 -294
rect 19929 68175 20239 76961
rect 21406 132594 21434 132599
rect 21406 74746 21434 132566
rect 28126 110138 28154 141526
rect 28182 124250 28210 142646
rect 28238 131306 28266 143206
rect 32224 137175 32384 137192
rect 32224 137147 32259 137175
rect 32287 137147 32321 137175
rect 32349 137147 32384 137175
rect 32224 137113 32384 137147
rect 32224 137085 32259 137113
rect 32287 137085 32321 137113
rect 32349 137085 32384 137113
rect 32224 137051 32384 137085
rect 32224 137023 32259 137051
rect 32287 137023 32321 137051
rect 32349 137023 32384 137051
rect 32224 136989 32384 137023
rect 32224 136961 32259 136989
rect 32287 136961 32321 136989
rect 32349 136961 32384 136989
rect 32224 136944 32384 136961
rect 33429 137175 33739 145961
rect 33429 137147 33477 137175
rect 33505 137147 33539 137175
rect 33567 137147 33601 137175
rect 33629 137147 33663 137175
rect 33691 137147 33739 137175
rect 33429 137113 33739 137147
rect 33429 137085 33477 137113
rect 33505 137085 33539 137113
rect 33567 137085 33601 137113
rect 33629 137085 33663 137113
rect 33691 137085 33739 137113
rect 33429 137051 33739 137085
rect 33429 137023 33477 137051
rect 33505 137023 33539 137051
rect 33567 137023 33601 137051
rect 33629 137023 33663 137051
rect 33691 137023 33739 137051
rect 33429 136989 33739 137023
rect 33429 136961 33477 136989
rect 33505 136961 33539 136989
rect 33567 136961 33601 136989
rect 33629 136961 33663 136989
rect 33691 136961 33739 136989
rect 28238 131273 28266 131278
rect 28182 124217 28210 124222
rect 33429 128175 33739 136961
rect 33429 128147 33477 128175
rect 33505 128147 33539 128175
rect 33567 128147 33601 128175
rect 33629 128147 33663 128175
rect 33691 128147 33739 128175
rect 33429 128113 33739 128147
rect 33429 128085 33477 128113
rect 33505 128085 33539 128113
rect 33567 128085 33601 128113
rect 33629 128085 33663 128113
rect 33691 128085 33739 128113
rect 33429 128051 33739 128085
rect 33429 128023 33477 128051
rect 33505 128023 33539 128051
rect 33567 128023 33601 128051
rect 33629 128023 33663 128051
rect 33691 128023 33739 128051
rect 33429 127989 33739 128023
rect 33429 127961 33477 127989
rect 33505 127961 33539 127989
rect 33567 127961 33601 127989
rect 33629 127961 33663 127989
rect 33691 127961 33739 127989
rect 28126 110105 28154 110110
rect 33429 119175 33739 127961
rect 33429 119147 33477 119175
rect 33505 119147 33539 119175
rect 33567 119147 33601 119175
rect 33629 119147 33663 119175
rect 33691 119147 33739 119175
rect 33429 119113 33739 119147
rect 33429 119085 33477 119113
rect 33505 119085 33539 119113
rect 33567 119085 33601 119113
rect 33629 119085 33663 119113
rect 33691 119085 33739 119113
rect 33429 119051 33739 119085
rect 33429 119023 33477 119051
rect 33505 119023 33539 119051
rect 33567 119023 33601 119051
rect 33629 119023 33663 119051
rect 33691 119023 33739 119051
rect 33429 118989 33739 119023
rect 33429 118961 33477 118989
rect 33505 118961 33539 118989
rect 33567 118961 33601 118989
rect 33629 118961 33663 118989
rect 33691 118961 33739 118989
rect 33429 110175 33739 118961
rect 33429 110147 33477 110175
rect 33505 110147 33539 110175
rect 33567 110147 33601 110175
rect 33629 110147 33663 110175
rect 33691 110147 33739 110175
rect 33429 110113 33739 110147
rect 33429 110085 33477 110113
rect 33505 110085 33539 110113
rect 33567 110085 33601 110113
rect 33629 110085 33663 110113
rect 33691 110085 33739 110113
rect 33429 110051 33739 110085
rect 33429 110023 33477 110051
rect 33505 110023 33539 110051
rect 33567 110023 33601 110051
rect 33629 110023 33663 110051
rect 33691 110023 33739 110051
rect 33429 109989 33739 110023
rect 33429 109961 33477 109989
rect 33505 109961 33539 109989
rect 33567 109961 33601 109989
rect 33629 109961 33663 109989
rect 33691 109961 33739 109989
rect 31584 101175 31744 101192
rect 31584 101147 31619 101175
rect 31647 101147 31681 101175
rect 31709 101147 31744 101175
rect 31584 101113 31744 101147
rect 31584 101085 31619 101113
rect 31647 101085 31681 101113
rect 31709 101085 31744 101113
rect 31584 101051 31744 101085
rect 31584 101023 31619 101051
rect 31647 101023 31681 101051
rect 31709 101023 31744 101051
rect 31584 100989 31744 101023
rect 31584 100961 31619 100989
rect 31647 100961 31681 100989
rect 31709 100961 31744 100989
rect 31584 100944 31744 100961
rect 33429 101175 33739 109961
rect 33429 101147 33477 101175
rect 33505 101147 33539 101175
rect 33567 101147 33601 101175
rect 33629 101147 33663 101175
rect 33691 101147 33739 101175
rect 33429 101113 33739 101147
rect 33429 101085 33477 101113
rect 33505 101085 33539 101113
rect 33567 101085 33601 101113
rect 33629 101085 33663 101113
rect 33691 101085 33739 101113
rect 33429 101051 33739 101085
rect 33429 101023 33477 101051
rect 33505 101023 33539 101051
rect 33567 101023 33601 101051
rect 33629 101023 33663 101051
rect 33691 101023 33739 101051
rect 33429 100989 33739 101023
rect 33429 100961 33477 100989
rect 33505 100961 33539 100989
rect 33567 100961 33601 100989
rect 33629 100961 33663 100989
rect 33691 100961 33739 100989
rect 23904 95175 24064 95192
rect 23904 95147 23939 95175
rect 23967 95147 24001 95175
rect 24029 95147 24064 95175
rect 23904 95113 24064 95147
rect 23904 95085 23939 95113
rect 23967 95085 24001 95113
rect 24029 95085 24064 95113
rect 23904 95051 24064 95085
rect 23904 95023 23939 95051
rect 23967 95023 24001 95051
rect 24029 95023 24064 95051
rect 23904 94989 24064 95023
rect 23904 94961 23939 94989
rect 23967 94961 24001 94989
rect 24029 94961 24064 94989
rect 23904 94944 24064 94961
rect 31584 92175 31744 92192
rect 31584 92147 31619 92175
rect 31647 92147 31681 92175
rect 31709 92147 31744 92175
rect 31584 92113 31744 92147
rect 31584 92085 31619 92113
rect 31647 92085 31681 92113
rect 31709 92085 31744 92113
rect 31584 92051 31744 92085
rect 31584 92023 31619 92051
rect 31647 92023 31681 92051
rect 31709 92023 31744 92051
rect 31584 91989 31744 92023
rect 31584 91961 31619 91989
rect 31647 91961 31681 91989
rect 31709 91961 31744 91989
rect 31584 91944 31744 91961
rect 33429 92175 33739 100961
rect 33429 92147 33477 92175
rect 33505 92147 33539 92175
rect 33567 92147 33601 92175
rect 33629 92147 33663 92175
rect 33691 92147 33739 92175
rect 33429 92113 33739 92147
rect 33429 92085 33477 92113
rect 33505 92085 33539 92113
rect 33567 92085 33601 92113
rect 33629 92085 33663 92113
rect 33691 92085 33739 92113
rect 33429 92051 33739 92085
rect 33429 92023 33477 92051
rect 33505 92023 33539 92051
rect 33567 92023 33601 92051
rect 33629 92023 33663 92051
rect 33691 92023 33739 92051
rect 33429 91989 33739 92023
rect 33429 91961 33477 91989
rect 33505 91961 33539 91989
rect 33567 91961 33601 91989
rect 33629 91961 33663 91989
rect 33691 91961 33739 91989
rect 33429 90103 33739 91961
rect 35289 167175 35599 170745
rect 35289 167147 35337 167175
rect 35365 167147 35399 167175
rect 35427 167147 35461 167175
rect 35489 167147 35523 167175
rect 35551 167147 35599 167175
rect 35289 167113 35599 167147
rect 35289 167085 35337 167113
rect 35365 167085 35399 167113
rect 35427 167085 35461 167113
rect 35489 167085 35523 167113
rect 35551 167085 35599 167113
rect 35289 167051 35599 167085
rect 35289 167023 35337 167051
rect 35365 167023 35399 167051
rect 35427 167023 35461 167051
rect 35489 167023 35523 167051
rect 35551 167023 35599 167051
rect 35289 166989 35599 167023
rect 35289 166961 35337 166989
rect 35365 166961 35399 166989
rect 35427 166961 35461 166989
rect 35489 166961 35523 166989
rect 35551 166961 35599 166989
rect 35289 158175 35599 166961
rect 48789 164175 49099 170745
rect 48789 164147 48837 164175
rect 48865 164147 48899 164175
rect 48927 164147 48961 164175
rect 48989 164147 49023 164175
rect 49051 164147 49099 164175
rect 48789 164113 49099 164147
rect 48789 164085 48837 164113
rect 48865 164085 48899 164113
rect 48927 164085 48961 164113
rect 48989 164085 49023 164113
rect 49051 164085 49099 164113
rect 48789 164051 49099 164085
rect 48789 164023 48837 164051
rect 48865 164023 48899 164051
rect 48927 164023 48961 164051
rect 48989 164023 49023 164051
rect 49051 164023 49099 164051
rect 48789 163989 49099 164023
rect 48789 163961 48837 163989
rect 48865 163961 48899 163989
rect 48927 163961 48961 163989
rect 48989 163961 49023 163989
rect 49051 163961 49099 163989
rect 35289 158147 35337 158175
rect 35365 158147 35399 158175
rect 35427 158147 35461 158175
rect 35489 158147 35523 158175
rect 35551 158147 35599 158175
rect 35289 158113 35599 158147
rect 35289 158085 35337 158113
rect 35365 158085 35399 158113
rect 35427 158085 35461 158113
rect 35489 158085 35523 158113
rect 35551 158085 35599 158113
rect 35289 158051 35599 158085
rect 35289 158023 35337 158051
rect 35365 158023 35399 158051
rect 35427 158023 35461 158051
rect 35489 158023 35523 158051
rect 35551 158023 35599 158051
rect 35289 157989 35599 158023
rect 35289 157961 35337 157989
rect 35365 157961 35399 157989
rect 35427 157961 35461 157989
rect 35489 157961 35523 157989
rect 35551 157961 35599 157989
rect 35289 149175 35599 157961
rect 39904 158175 40064 158192
rect 39904 158147 39939 158175
rect 39967 158147 40001 158175
rect 40029 158147 40064 158175
rect 39904 158113 40064 158147
rect 39904 158085 39939 158113
rect 39967 158085 40001 158113
rect 40029 158085 40064 158113
rect 39904 158051 40064 158085
rect 39904 158023 39939 158051
rect 39967 158023 40001 158051
rect 40029 158023 40064 158051
rect 39904 157989 40064 158023
rect 39904 157961 39939 157989
rect 39967 157961 40001 157989
rect 40029 157961 40064 157989
rect 39904 157944 40064 157961
rect 47584 155175 47744 155192
rect 47584 155147 47619 155175
rect 47647 155147 47681 155175
rect 47709 155147 47744 155175
rect 47584 155113 47744 155147
rect 47584 155085 47619 155113
rect 47647 155085 47681 155113
rect 47709 155085 47744 155113
rect 47584 155051 47744 155085
rect 47584 155023 47619 155051
rect 47647 155023 47681 155051
rect 47709 155023 47744 155051
rect 47584 154989 47744 155023
rect 47584 154961 47619 154989
rect 47647 154961 47681 154989
rect 47709 154961 47744 154989
rect 47584 154944 47744 154961
rect 48789 155175 49099 163961
rect 48789 155147 48837 155175
rect 48865 155147 48899 155175
rect 48927 155147 48961 155175
rect 48989 155147 49023 155175
rect 49051 155147 49099 155175
rect 48789 155113 49099 155147
rect 48789 155085 48837 155113
rect 48865 155085 48899 155113
rect 48927 155085 48961 155113
rect 48989 155085 49023 155113
rect 49051 155085 49099 155113
rect 48789 155051 49099 155085
rect 48789 155023 48837 155051
rect 48865 155023 48899 155051
rect 48927 155023 48961 155051
rect 48989 155023 49023 155051
rect 49051 155023 49099 155051
rect 48789 154989 49099 155023
rect 48789 154961 48837 154989
rect 48865 154961 48899 154989
rect 48927 154961 48961 154989
rect 48989 154961 49023 154989
rect 49051 154961 49099 154989
rect 35289 149147 35337 149175
rect 35365 149147 35399 149175
rect 35427 149147 35461 149175
rect 35489 149147 35523 149175
rect 35551 149147 35599 149175
rect 35289 149113 35599 149147
rect 35289 149085 35337 149113
rect 35365 149085 35399 149113
rect 35427 149085 35461 149113
rect 35489 149085 35523 149113
rect 35551 149085 35599 149113
rect 35289 149051 35599 149085
rect 35289 149023 35337 149051
rect 35365 149023 35399 149051
rect 35427 149023 35461 149051
rect 35489 149023 35523 149051
rect 35551 149023 35599 149051
rect 35289 148989 35599 149023
rect 35289 148961 35337 148989
rect 35365 148961 35399 148989
rect 35427 148961 35461 148989
rect 35489 148961 35523 148989
rect 35551 148961 35599 148989
rect 35289 140175 35599 148961
rect 39904 149175 40064 149192
rect 39904 149147 39939 149175
rect 39967 149147 40001 149175
rect 40029 149147 40064 149175
rect 39904 149113 40064 149147
rect 39904 149085 39939 149113
rect 39967 149085 40001 149113
rect 40029 149085 40064 149113
rect 39904 149051 40064 149085
rect 39904 149023 39939 149051
rect 39967 149023 40001 149051
rect 40029 149023 40064 149051
rect 39904 148989 40064 149023
rect 39904 148961 39939 148989
rect 39967 148961 40001 148989
rect 40029 148961 40064 148989
rect 39904 148944 40064 148961
rect 47584 146175 47744 146192
rect 47584 146147 47619 146175
rect 47647 146147 47681 146175
rect 47709 146147 47744 146175
rect 47584 146113 47744 146147
rect 47584 146085 47619 146113
rect 47647 146085 47681 146113
rect 47709 146085 47744 146113
rect 47584 146051 47744 146085
rect 47584 146023 47619 146051
rect 47647 146023 47681 146051
rect 47709 146023 47744 146051
rect 47584 145989 47744 146023
rect 47584 145961 47619 145989
rect 47647 145961 47681 145989
rect 47709 145961 47744 145989
rect 47584 145944 47744 145961
rect 48789 146175 49099 154961
rect 48789 146147 48837 146175
rect 48865 146147 48899 146175
rect 48927 146147 48961 146175
rect 48989 146147 49023 146175
rect 49051 146147 49099 146175
rect 48789 146113 49099 146147
rect 48789 146085 48837 146113
rect 48865 146085 48899 146113
rect 48927 146085 48961 146113
rect 48989 146085 49023 146113
rect 49051 146085 49099 146113
rect 48789 146051 49099 146085
rect 48789 146023 48837 146051
rect 48865 146023 48899 146051
rect 48927 146023 48961 146051
rect 48989 146023 49023 146051
rect 49051 146023 49099 146051
rect 48789 145989 49099 146023
rect 48789 145961 48837 145989
rect 48865 145961 48899 145989
rect 48927 145961 48961 145989
rect 48989 145961 49023 145989
rect 49051 145961 49099 145989
rect 35289 140147 35337 140175
rect 35365 140147 35399 140175
rect 35427 140147 35461 140175
rect 35489 140147 35523 140175
rect 35551 140147 35599 140175
rect 35289 140113 35599 140147
rect 35289 140085 35337 140113
rect 35365 140085 35399 140113
rect 35427 140085 35461 140113
rect 35489 140085 35523 140113
rect 35551 140085 35599 140113
rect 35289 140051 35599 140085
rect 35289 140023 35337 140051
rect 35365 140023 35399 140051
rect 35427 140023 35461 140051
rect 35489 140023 35523 140051
rect 35551 140023 35599 140051
rect 35289 139989 35599 140023
rect 35289 139961 35337 139989
rect 35365 139961 35399 139989
rect 35427 139961 35461 139989
rect 35489 139961 35523 139989
rect 35551 139961 35599 139989
rect 35289 131175 35599 139961
rect 39904 140175 40064 140192
rect 39904 140147 39939 140175
rect 39967 140147 40001 140175
rect 40029 140147 40064 140175
rect 39904 140113 40064 140147
rect 39904 140085 39939 140113
rect 39967 140085 40001 140113
rect 40029 140085 40064 140113
rect 39904 140051 40064 140085
rect 39904 140023 39939 140051
rect 39967 140023 40001 140051
rect 40029 140023 40064 140051
rect 39904 139989 40064 140023
rect 39904 139961 39939 139989
rect 39967 139961 40001 139989
rect 40029 139961 40064 139989
rect 39904 139944 40064 139961
rect 47584 137175 47744 137192
rect 47584 137147 47619 137175
rect 47647 137147 47681 137175
rect 47709 137147 47744 137175
rect 47584 137113 47744 137147
rect 47584 137085 47619 137113
rect 47647 137085 47681 137113
rect 47709 137085 47744 137113
rect 47584 137051 47744 137085
rect 47584 137023 47619 137051
rect 47647 137023 47681 137051
rect 47709 137023 47744 137051
rect 47584 136989 47744 137023
rect 47584 136961 47619 136989
rect 47647 136961 47681 136989
rect 47709 136961 47744 136989
rect 47584 136944 47744 136961
rect 48789 137175 49099 145961
rect 48789 137147 48837 137175
rect 48865 137147 48899 137175
rect 48927 137147 48961 137175
rect 48989 137147 49023 137175
rect 49051 137147 49099 137175
rect 48789 137113 49099 137147
rect 48789 137085 48837 137113
rect 48865 137085 48899 137113
rect 48927 137085 48961 137113
rect 48989 137085 49023 137113
rect 49051 137085 49099 137113
rect 48789 137051 49099 137085
rect 48789 137023 48837 137051
rect 48865 137023 48899 137051
rect 48927 137023 48961 137051
rect 48989 137023 49023 137051
rect 49051 137023 49099 137051
rect 48789 136989 49099 137023
rect 48789 136961 48837 136989
rect 48865 136961 48899 136989
rect 48927 136961 48961 136989
rect 48989 136961 49023 136989
rect 49051 136961 49099 136989
rect 35289 131147 35337 131175
rect 35365 131147 35399 131175
rect 35427 131147 35461 131175
rect 35489 131147 35523 131175
rect 35551 131147 35599 131175
rect 35289 131113 35599 131147
rect 35289 131085 35337 131113
rect 35365 131085 35399 131113
rect 35427 131085 35461 131113
rect 35489 131085 35523 131113
rect 35551 131085 35599 131113
rect 35289 131051 35599 131085
rect 35289 131023 35337 131051
rect 35365 131023 35399 131051
rect 35427 131023 35461 131051
rect 35489 131023 35523 131051
rect 35551 131023 35599 131051
rect 35289 130989 35599 131023
rect 35289 130961 35337 130989
rect 35365 130961 35399 130989
rect 35427 130961 35461 130989
rect 35489 130961 35523 130989
rect 35551 130961 35599 130989
rect 35289 122175 35599 130961
rect 35289 122147 35337 122175
rect 35365 122147 35399 122175
rect 35427 122147 35461 122175
rect 35489 122147 35523 122175
rect 35551 122147 35599 122175
rect 35289 122113 35599 122147
rect 35289 122085 35337 122113
rect 35365 122085 35399 122113
rect 35427 122085 35461 122113
rect 35489 122085 35523 122113
rect 35551 122085 35599 122113
rect 35289 122051 35599 122085
rect 35289 122023 35337 122051
rect 35365 122023 35399 122051
rect 35427 122023 35461 122051
rect 35489 122023 35523 122051
rect 35551 122023 35599 122051
rect 35289 121989 35599 122023
rect 35289 121961 35337 121989
rect 35365 121961 35399 121989
rect 35427 121961 35461 121989
rect 35489 121961 35523 121989
rect 35551 121961 35599 121989
rect 35289 113175 35599 121961
rect 35289 113147 35337 113175
rect 35365 113147 35399 113175
rect 35427 113147 35461 113175
rect 35489 113147 35523 113175
rect 35551 113147 35599 113175
rect 35289 113113 35599 113147
rect 35289 113085 35337 113113
rect 35365 113085 35399 113113
rect 35427 113085 35461 113113
rect 35489 113085 35523 113113
rect 35551 113085 35599 113113
rect 35289 113051 35599 113085
rect 35289 113023 35337 113051
rect 35365 113023 35399 113051
rect 35427 113023 35461 113051
rect 35489 113023 35523 113051
rect 35551 113023 35599 113051
rect 35289 112989 35599 113023
rect 35289 112961 35337 112989
rect 35365 112961 35399 112989
rect 35427 112961 35461 112989
rect 35489 112961 35523 112989
rect 35551 112961 35599 112989
rect 35289 104175 35599 112961
rect 35289 104147 35337 104175
rect 35365 104147 35399 104175
rect 35427 104147 35461 104175
rect 35489 104147 35523 104175
rect 35551 104147 35599 104175
rect 35289 104113 35599 104147
rect 35289 104085 35337 104113
rect 35365 104085 35399 104113
rect 35427 104085 35461 104113
rect 35489 104085 35523 104113
rect 35551 104085 35599 104113
rect 35289 104051 35599 104085
rect 35289 104023 35337 104051
rect 35365 104023 35399 104051
rect 35427 104023 35461 104051
rect 35489 104023 35523 104051
rect 35551 104023 35599 104051
rect 35289 103989 35599 104023
rect 35289 103961 35337 103989
rect 35365 103961 35399 103989
rect 35427 103961 35461 103989
rect 35489 103961 35523 103989
rect 35551 103961 35599 103989
rect 35289 95175 35599 103961
rect 48789 128175 49099 136961
rect 48789 128147 48837 128175
rect 48865 128147 48899 128175
rect 48927 128147 48961 128175
rect 48989 128147 49023 128175
rect 49051 128147 49099 128175
rect 48789 128113 49099 128147
rect 48789 128085 48837 128113
rect 48865 128085 48899 128113
rect 48927 128085 48961 128113
rect 48989 128085 49023 128113
rect 49051 128085 49099 128113
rect 48789 128051 49099 128085
rect 48789 128023 48837 128051
rect 48865 128023 48899 128051
rect 48927 128023 48961 128051
rect 48989 128023 49023 128051
rect 49051 128023 49099 128051
rect 48789 127989 49099 128023
rect 48789 127961 48837 127989
rect 48865 127961 48899 127989
rect 48927 127961 48961 127989
rect 48989 127961 49023 127989
rect 49051 127961 49099 127989
rect 48789 119175 49099 127961
rect 48789 119147 48837 119175
rect 48865 119147 48899 119175
rect 48927 119147 48961 119175
rect 48989 119147 49023 119175
rect 49051 119147 49099 119175
rect 48789 119113 49099 119147
rect 48789 119085 48837 119113
rect 48865 119085 48899 119113
rect 48927 119085 48961 119113
rect 48989 119085 49023 119113
rect 49051 119085 49099 119113
rect 48789 119051 49099 119085
rect 48789 119023 48837 119051
rect 48865 119023 48899 119051
rect 48927 119023 48961 119051
rect 48989 119023 49023 119051
rect 49051 119023 49099 119051
rect 48789 118989 49099 119023
rect 48789 118961 48837 118989
rect 48865 118961 48899 118989
rect 48927 118961 48961 118989
rect 48989 118961 49023 118989
rect 49051 118961 49099 118989
rect 48789 110175 49099 118961
rect 48789 110147 48837 110175
rect 48865 110147 48899 110175
rect 48927 110147 48961 110175
rect 48989 110147 49023 110175
rect 49051 110147 49099 110175
rect 48789 110113 49099 110147
rect 48789 110085 48837 110113
rect 48865 110085 48899 110113
rect 48927 110085 48961 110113
rect 48989 110085 49023 110113
rect 49051 110085 49099 110113
rect 48789 110051 49099 110085
rect 48789 110023 48837 110051
rect 48865 110023 48899 110051
rect 48927 110023 48961 110051
rect 48989 110023 49023 110051
rect 49051 110023 49099 110051
rect 48789 109989 49099 110023
rect 48789 109961 48837 109989
rect 48865 109961 48899 109989
rect 48927 109961 48961 109989
rect 48989 109961 49023 109989
rect 49051 109961 49099 109989
rect 46944 101175 47104 101192
rect 46944 101147 46979 101175
rect 47007 101147 47041 101175
rect 47069 101147 47104 101175
rect 46944 101113 47104 101147
rect 46944 101085 46979 101113
rect 47007 101085 47041 101113
rect 47069 101085 47104 101113
rect 46944 101051 47104 101085
rect 46944 101023 46979 101051
rect 47007 101023 47041 101051
rect 47069 101023 47104 101051
rect 46944 100989 47104 101023
rect 46944 100961 46979 100989
rect 47007 100961 47041 100989
rect 47069 100961 47104 100989
rect 46944 100944 47104 100961
rect 48789 101175 49099 109961
rect 48789 101147 48837 101175
rect 48865 101147 48899 101175
rect 48927 101147 48961 101175
rect 48989 101147 49023 101175
rect 49051 101147 49099 101175
rect 48789 101113 49099 101147
rect 48789 101085 48837 101113
rect 48865 101085 48899 101113
rect 48927 101085 48961 101113
rect 48989 101085 49023 101113
rect 49051 101085 49099 101113
rect 48789 101051 49099 101085
rect 48789 101023 48837 101051
rect 48865 101023 48899 101051
rect 48927 101023 48961 101051
rect 48989 101023 49023 101051
rect 49051 101023 49099 101051
rect 48789 100989 49099 101023
rect 48789 100961 48837 100989
rect 48865 100961 48899 100989
rect 48927 100961 48961 100989
rect 48989 100961 49023 100989
rect 49051 100961 49099 100989
rect 35289 95147 35337 95175
rect 35365 95147 35399 95175
rect 35427 95147 35461 95175
rect 35489 95147 35523 95175
rect 35551 95147 35599 95175
rect 35289 95113 35599 95147
rect 35289 95085 35337 95113
rect 35365 95085 35399 95113
rect 35427 95085 35461 95113
rect 35489 95085 35523 95113
rect 35551 95085 35599 95113
rect 35289 95051 35599 95085
rect 35289 95023 35337 95051
rect 35365 95023 35399 95051
rect 35427 95023 35461 95051
rect 35489 95023 35523 95051
rect 35551 95023 35599 95051
rect 35289 94989 35599 95023
rect 35289 94961 35337 94989
rect 35365 94961 35399 94989
rect 35427 94961 35461 94989
rect 35489 94961 35523 94989
rect 35551 94961 35599 94989
rect 35289 90103 35599 94961
rect 39264 95175 39424 95192
rect 39264 95147 39299 95175
rect 39327 95147 39361 95175
rect 39389 95147 39424 95175
rect 39264 95113 39424 95147
rect 39264 95085 39299 95113
rect 39327 95085 39361 95113
rect 39389 95085 39424 95113
rect 39264 95051 39424 95085
rect 39264 95023 39299 95051
rect 39327 95023 39361 95051
rect 39389 95023 39424 95051
rect 39264 94989 39424 95023
rect 39264 94961 39299 94989
rect 39327 94961 39361 94989
rect 39389 94961 39424 94989
rect 39264 94944 39424 94961
rect 46944 92175 47104 92192
rect 46944 92147 46979 92175
rect 47007 92147 47041 92175
rect 47069 92147 47104 92175
rect 46944 92113 47104 92147
rect 46944 92085 46979 92113
rect 47007 92085 47041 92113
rect 47069 92085 47104 92113
rect 46944 92051 47104 92085
rect 46944 92023 46979 92051
rect 47007 92023 47041 92051
rect 47069 92023 47104 92051
rect 46944 91989 47104 92023
rect 46944 91961 46979 91989
rect 47007 91961 47041 91989
rect 47069 91961 47104 91989
rect 46944 91944 47104 91961
rect 48789 92175 49099 100961
rect 48789 92147 48837 92175
rect 48865 92147 48899 92175
rect 48927 92147 48961 92175
rect 48989 92147 49023 92175
rect 49051 92147 49099 92175
rect 48789 92113 49099 92147
rect 48789 92085 48837 92113
rect 48865 92085 48899 92113
rect 48927 92085 48961 92113
rect 48989 92085 49023 92113
rect 49051 92085 49099 92113
rect 48789 92051 49099 92085
rect 48789 92023 48837 92051
rect 48865 92023 48899 92051
rect 48927 92023 48961 92051
rect 48989 92023 49023 92051
rect 49051 92023 49099 92051
rect 48789 91989 49099 92023
rect 48789 91961 48837 91989
rect 48865 91961 48899 91989
rect 48927 91961 48961 91989
rect 48989 91961 49023 91989
rect 49051 91961 49099 91989
rect 48789 90103 49099 91961
rect 50649 167175 50959 170745
rect 50649 167147 50697 167175
rect 50725 167147 50759 167175
rect 50787 167147 50821 167175
rect 50849 167147 50883 167175
rect 50911 167147 50959 167175
rect 50649 167113 50959 167147
rect 50649 167085 50697 167113
rect 50725 167085 50759 167113
rect 50787 167085 50821 167113
rect 50849 167085 50883 167113
rect 50911 167085 50959 167113
rect 50649 167051 50959 167085
rect 50649 167023 50697 167051
rect 50725 167023 50759 167051
rect 50787 167023 50821 167051
rect 50849 167023 50883 167051
rect 50911 167023 50959 167051
rect 50649 166989 50959 167023
rect 50649 166961 50697 166989
rect 50725 166961 50759 166989
rect 50787 166961 50821 166989
rect 50849 166961 50883 166989
rect 50911 166961 50959 166989
rect 50649 158175 50959 166961
rect 64149 164175 64459 170745
rect 64149 164147 64197 164175
rect 64225 164147 64259 164175
rect 64287 164147 64321 164175
rect 64349 164147 64383 164175
rect 64411 164147 64459 164175
rect 64149 164113 64459 164147
rect 64149 164085 64197 164113
rect 64225 164085 64259 164113
rect 64287 164085 64321 164113
rect 64349 164085 64383 164113
rect 64411 164085 64459 164113
rect 64149 164051 64459 164085
rect 64149 164023 64197 164051
rect 64225 164023 64259 164051
rect 64287 164023 64321 164051
rect 64349 164023 64383 164051
rect 64411 164023 64459 164051
rect 64149 163989 64459 164023
rect 64149 163961 64197 163989
rect 64225 163961 64259 163989
rect 64287 163961 64321 163989
rect 64349 163961 64383 163989
rect 64411 163961 64459 163989
rect 50649 158147 50697 158175
rect 50725 158147 50759 158175
rect 50787 158147 50821 158175
rect 50849 158147 50883 158175
rect 50911 158147 50959 158175
rect 50649 158113 50959 158147
rect 50649 158085 50697 158113
rect 50725 158085 50759 158113
rect 50787 158085 50821 158113
rect 50849 158085 50883 158113
rect 50911 158085 50959 158113
rect 50649 158051 50959 158085
rect 50649 158023 50697 158051
rect 50725 158023 50759 158051
rect 50787 158023 50821 158051
rect 50849 158023 50883 158051
rect 50911 158023 50959 158051
rect 50649 157989 50959 158023
rect 50649 157961 50697 157989
rect 50725 157961 50759 157989
rect 50787 157961 50821 157989
rect 50849 157961 50883 157989
rect 50911 157961 50959 157989
rect 50649 149175 50959 157961
rect 55264 158175 55424 158192
rect 55264 158147 55299 158175
rect 55327 158147 55361 158175
rect 55389 158147 55424 158175
rect 55264 158113 55424 158147
rect 55264 158085 55299 158113
rect 55327 158085 55361 158113
rect 55389 158085 55424 158113
rect 55264 158051 55424 158085
rect 55264 158023 55299 158051
rect 55327 158023 55361 158051
rect 55389 158023 55424 158051
rect 55264 157989 55424 158023
rect 55264 157961 55299 157989
rect 55327 157961 55361 157989
rect 55389 157961 55424 157989
rect 55264 157944 55424 157961
rect 62944 155175 63104 155192
rect 62944 155147 62979 155175
rect 63007 155147 63041 155175
rect 63069 155147 63104 155175
rect 62944 155113 63104 155147
rect 62944 155085 62979 155113
rect 63007 155085 63041 155113
rect 63069 155085 63104 155113
rect 62944 155051 63104 155085
rect 62944 155023 62979 155051
rect 63007 155023 63041 155051
rect 63069 155023 63104 155051
rect 62944 154989 63104 155023
rect 62944 154961 62979 154989
rect 63007 154961 63041 154989
rect 63069 154961 63104 154989
rect 62944 154944 63104 154961
rect 64149 155175 64459 163961
rect 64149 155147 64197 155175
rect 64225 155147 64259 155175
rect 64287 155147 64321 155175
rect 64349 155147 64383 155175
rect 64411 155147 64459 155175
rect 64149 155113 64459 155147
rect 64149 155085 64197 155113
rect 64225 155085 64259 155113
rect 64287 155085 64321 155113
rect 64349 155085 64383 155113
rect 64411 155085 64459 155113
rect 64149 155051 64459 155085
rect 64149 155023 64197 155051
rect 64225 155023 64259 155051
rect 64287 155023 64321 155051
rect 64349 155023 64383 155051
rect 64411 155023 64459 155051
rect 64149 154989 64459 155023
rect 64149 154961 64197 154989
rect 64225 154961 64259 154989
rect 64287 154961 64321 154989
rect 64349 154961 64383 154989
rect 64411 154961 64459 154989
rect 50649 149147 50697 149175
rect 50725 149147 50759 149175
rect 50787 149147 50821 149175
rect 50849 149147 50883 149175
rect 50911 149147 50959 149175
rect 50649 149113 50959 149147
rect 50649 149085 50697 149113
rect 50725 149085 50759 149113
rect 50787 149085 50821 149113
rect 50849 149085 50883 149113
rect 50911 149085 50959 149113
rect 50649 149051 50959 149085
rect 50649 149023 50697 149051
rect 50725 149023 50759 149051
rect 50787 149023 50821 149051
rect 50849 149023 50883 149051
rect 50911 149023 50959 149051
rect 50649 148989 50959 149023
rect 50649 148961 50697 148989
rect 50725 148961 50759 148989
rect 50787 148961 50821 148989
rect 50849 148961 50883 148989
rect 50911 148961 50959 148989
rect 50649 140175 50959 148961
rect 55264 149175 55424 149192
rect 55264 149147 55299 149175
rect 55327 149147 55361 149175
rect 55389 149147 55424 149175
rect 55264 149113 55424 149147
rect 55264 149085 55299 149113
rect 55327 149085 55361 149113
rect 55389 149085 55424 149113
rect 55264 149051 55424 149085
rect 55264 149023 55299 149051
rect 55327 149023 55361 149051
rect 55389 149023 55424 149051
rect 55264 148989 55424 149023
rect 55264 148961 55299 148989
rect 55327 148961 55361 148989
rect 55389 148961 55424 148989
rect 55264 148944 55424 148961
rect 62944 146175 63104 146192
rect 62944 146147 62979 146175
rect 63007 146147 63041 146175
rect 63069 146147 63104 146175
rect 62944 146113 63104 146147
rect 62944 146085 62979 146113
rect 63007 146085 63041 146113
rect 63069 146085 63104 146113
rect 62944 146051 63104 146085
rect 62944 146023 62979 146051
rect 63007 146023 63041 146051
rect 63069 146023 63104 146051
rect 62944 145989 63104 146023
rect 62944 145961 62979 145989
rect 63007 145961 63041 145989
rect 63069 145961 63104 145989
rect 62944 145944 63104 145961
rect 64149 146175 64459 154961
rect 64149 146147 64197 146175
rect 64225 146147 64259 146175
rect 64287 146147 64321 146175
rect 64349 146147 64383 146175
rect 64411 146147 64459 146175
rect 64149 146113 64459 146147
rect 64149 146085 64197 146113
rect 64225 146085 64259 146113
rect 64287 146085 64321 146113
rect 64349 146085 64383 146113
rect 64411 146085 64459 146113
rect 64149 146051 64459 146085
rect 64149 146023 64197 146051
rect 64225 146023 64259 146051
rect 64287 146023 64321 146051
rect 64349 146023 64383 146051
rect 64411 146023 64459 146051
rect 64149 145989 64459 146023
rect 64149 145961 64197 145989
rect 64225 145961 64259 145989
rect 64287 145961 64321 145989
rect 64349 145961 64383 145989
rect 64411 145961 64459 145989
rect 50649 140147 50697 140175
rect 50725 140147 50759 140175
rect 50787 140147 50821 140175
rect 50849 140147 50883 140175
rect 50911 140147 50959 140175
rect 50649 140113 50959 140147
rect 50649 140085 50697 140113
rect 50725 140085 50759 140113
rect 50787 140085 50821 140113
rect 50849 140085 50883 140113
rect 50911 140085 50959 140113
rect 50649 140051 50959 140085
rect 50649 140023 50697 140051
rect 50725 140023 50759 140051
rect 50787 140023 50821 140051
rect 50849 140023 50883 140051
rect 50911 140023 50959 140051
rect 50649 139989 50959 140023
rect 50649 139961 50697 139989
rect 50725 139961 50759 139989
rect 50787 139961 50821 139989
rect 50849 139961 50883 139989
rect 50911 139961 50959 139989
rect 50649 131175 50959 139961
rect 55264 140175 55424 140192
rect 55264 140147 55299 140175
rect 55327 140147 55361 140175
rect 55389 140147 55424 140175
rect 55264 140113 55424 140147
rect 55264 140085 55299 140113
rect 55327 140085 55361 140113
rect 55389 140085 55424 140113
rect 55264 140051 55424 140085
rect 55264 140023 55299 140051
rect 55327 140023 55361 140051
rect 55389 140023 55424 140051
rect 55264 139989 55424 140023
rect 55264 139961 55299 139989
rect 55327 139961 55361 139989
rect 55389 139961 55424 139989
rect 55264 139944 55424 139961
rect 62944 137175 63104 137192
rect 62944 137147 62979 137175
rect 63007 137147 63041 137175
rect 63069 137147 63104 137175
rect 62944 137113 63104 137147
rect 62944 137085 62979 137113
rect 63007 137085 63041 137113
rect 63069 137085 63104 137113
rect 62944 137051 63104 137085
rect 62944 137023 62979 137051
rect 63007 137023 63041 137051
rect 63069 137023 63104 137051
rect 62944 136989 63104 137023
rect 62944 136961 62979 136989
rect 63007 136961 63041 136989
rect 63069 136961 63104 136989
rect 62944 136944 63104 136961
rect 64149 137175 64459 145961
rect 64149 137147 64197 137175
rect 64225 137147 64259 137175
rect 64287 137147 64321 137175
rect 64349 137147 64383 137175
rect 64411 137147 64459 137175
rect 64149 137113 64459 137147
rect 64149 137085 64197 137113
rect 64225 137085 64259 137113
rect 64287 137085 64321 137113
rect 64349 137085 64383 137113
rect 64411 137085 64459 137113
rect 64149 137051 64459 137085
rect 64149 137023 64197 137051
rect 64225 137023 64259 137051
rect 64287 137023 64321 137051
rect 64349 137023 64383 137051
rect 64411 137023 64459 137051
rect 64149 136989 64459 137023
rect 64149 136961 64197 136989
rect 64225 136961 64259 136989
rect 64287 136961 64321 136989
rect 64349 136961 64383 136989
rect 64411 136961 64459 136989
rect 50649 131147 50697 131175
rect 50725 131147 50759 131175
rect 50787 131147 50821 131175
rect 50849 131147 50883 131175
rect 50911 131147 50959 131175
rect 50649 131113 50959 131147
rect 50649 131085 50697 131113
rect 50725 131085 50759 131113
rect 50787 131085 50821 131113
rect 50849 131085 50883 131113
rect 50911 131085 50959 131113
rect 50649 131051 50959 131085
rect 50649 131023 50697 131051
rect 50725 131023 50759 131051
rect 50787 131023 50821 131051
rect 50849 131023 50883 131051
rect 50911 131023 50959 131051
rect 50649 130989 50959 131023
rect 50649 130961 50697 130989
rect 50725 130961 50759 130989
rect 50787 130961 50821 130989
rect 50849 130961 50883 130989
rect 50911 130961 50959 130989
rect 50649 122175 50959 130961
rect 50649 122147 50697 122175
rect 50725 122147 50759 122175
rect 50787 122147 50821 122175
rect 50849 122147 50883 122175
rect 50911 122147 50959 122175
rect 50649 122113 50959 122147
rect 50649 122085 50697 122113
rect 50725 122085 50759 122113
rect 50787 122085 50821 122113
rect 50849 122085 50883 122113
rect 50911 122085 50959 122113
rect 50649 122051 50959 122085
rect 50649 122023 50697 122051
rect 50725 122023 50759 122051
rect 50787 122023 50821 122051
rect 50849 122023 50883 122051
rect 50911 122023 50959 122051
rect 50649 121989 50959 122023
rect 50649 121961 50697 121989
rect 50725 121961 50759 121989
rect 50787 121961 50821 121989
rect 50849 121961 50883 121989
rect 50911 121961 50959 121989
rect 50649 113175 50959 121961
rect 50649 113147 50697 113175
rect 50725 113147 50759 113175
rect 50787 113147 50821 113175
rect 50849 113147 50883 113175
rect 50911 113147 50959 113175
rect 50649 113113 50959 113147
rect 50649 113085 50697 113113
rect 50725 113085 50759 113113
rect 50787 113085 50821 113113
rect 50849 113085 50883 113113
rect 50911 113085 50959 113113
rect 50649 113051 50959 113085
rect 50649 113023 50697 113051
rect 50725 113023 50759 113051
rect 50787 113023 50821 113051
rect 50849 113023 50883 113051
rect 50911 113023 50959 113051
rect 50649 112989 50959 113023
rect 50649 112961 50697 112989
rect 50725 112961 50759 112989
rect 50787 112961 50821 112989
rect 50849 112961 50883 112989
rect 50911 112961 50959 112989
rect 50649 104175 50959 112961
rect 50649 104147 50697 104175
rect 50725 104147 50759 104175
rect 50787 104147 50821 104175
rect 50849 104147 50883 104175
rect 50911 104147 50959 104175
rect 50649 104113 50959 104147
rect 50649 104085 50697 104113
rect 50725 104085 50759 104113
rect 50787 104085 50821 104113
rect 50849 104085 50883 104113
rect 50911 104085 50959 104113
rect 50649 104051 50959 104085
rect 50649 104023 50697 104051
rect 50725 104023 50759 104051
rect 50787 104023 50821 104051
rect 50849 104023 50883 104051
rect 50911 104023 50959 104051
rect 50649 103989 50959 104023
rect 50649 103961 50697 103989
rect 50725 103961 50759 103989
rect 50787 103961 50821 103989
rect 50849 103961 50883 103989
rect 50911 103961 50959 103989
rect 50649 95175 50959 103961
rect 64149 128175 64459 136961
rect 64149 128147 64197 128175
rect 64225 128147 64259 128175
rect 64287 128147 64321 128175
rect 64349 128147 64383 128175
rect 64411 128147 64459 128175
rect 64149 128113 64459 128147
rect 64149 128085 64197 128113
rect 64225 128085 64259 128113
rect 64287 128085 64321 128113
rect 64349 128085 64383 128113
rect 64411 128085 64459 128113
rect 64149 128051 64459 128085
rect 64149 128023 64197 128051
rect 64225 128023 64259 128051
rect 64287 128023 64321 128051
rect 64349 128023 64383 128051
rect 64411 128023 64459 128051
rect 64149 127989 64459 128023
rect 64149 127961 64197 127989
rect 64225 127961 64259 127989
rect 64287 127961 64321 127989
rect 64349 127961 64383 127989
rect 64411 127961 64459 127989
rect 64149 119175 64459 127961
rect 64149 119147 64197 119175
rect 64225 119147 64259 119175
rect 64287 119147 64321 119175
rect 64349 119147 64383 119175
rect 64411 119147 64459 119175
rect 64149 119113 64459 119147
rect 64149 119085 64197 119113
rect 64225 119085 64259 119113
rect 64287 119085 64321 119113
rect 64349 119085 64383 119113
rect 64411 119085 64459 119113
rect 64149 119051 64459 119085
rect 64149 119023 64197 119051
rect 64225 119023 64259 119051
rect 64287 119023 64321 119051
rect 64349 119023 64383 119051
rect 64411 119023 64459 119051
rect 64149 118989 64459 119023
rect 64149 118961 64197 118989
rect 64225 118961 64259 118989
rect 64287 118961 64321 118989
rect 64349 118961 64383 118989
rect 64411 118961 64459 118989
rect 64149 110175 64459 118961
rect 64149 110147 64197 110175
rect 64225 110147 64259 110175
rect 64287 110147 64321 110175
rect 64349 110147 64383 110175
rect 64411 110147 64459 110175
rect 64149 110113 64459 110147
rect 64149 110085 64197 110113
rect 64225 110085 64259 110113
rect 64287 110085 64321 110113
rect 64349 110085 64383 110113
rect 64411 110085 64459 110113
rect 64149 110051 64459 110085
rect 64149 110023 64197 110051
rect 64225 110023 64259 110051
rect 64287 110023 64321 110051
rect 64349 110023 64383 110051
rect 64411 110023 64459 110051
rect 64149 109989 64459 110023
rect 64149 109961 64197 109989
rect 64225 109961 64259 109989
rect 64287 109961 64321 109989
rect 64349 109961 64383 109989
rect 64411 109961 64459 109989
rect 62304 101175 62464 101192
rect 62304 101147 62339 101175
rect 62367 101147 62401 101175
rect 62429 101147 62464 101175
rect 62304 101113 62464 101147
rect 62304 101085 62339 101113
rect 62367 101085 62401 101113
rect 62429 101085 62464 101113
rect 62304 101051 62464 101085
rect 62304 101023 62339 101051
rect 62367 101023 62401 101051
rect 62429 101023 62464 101051
rect 62304 100989 62464 101023
rect 62304 100961 62339 100989
rect 62367 100961 62401 100989
rect 62429 100961 62464 100989
rect 62304 100944 62464 100961
rect 64149 101175 64459 109961
rect 64149 101147 64197 101175
rect 64225 101147 64259 101175
rect 64287 101147 64321 101175
rect 64349 101147 64383 101175
rect 64411 101147 64459 101175
rect 64149 101113 64459 101147
rect 64149 101085 64197 101113
rect 64225 101085 64259 101113
rect 64287 101085 64321 101113
rect 64349 101085 64383 101113
rect 64411 101085 64459 101113
rect 64149 101051 64459 101085
rect 64149 101023 64197 101051
rect 64225 101023 64259 101051
rect 64287 101023 64321 101051
rect 64349 101023 64383 101051
rect 64411 101023 64459 101051
rect 64149 100989 64459 101023
rect 64149 100961 64197 100989
rect 64225 100961 64259 100989
rect 64287 100961 64321 100989
rect 64349 100961 64383 100989
rect 64411 100961 64459 100989
rect 50649 95147 50697 95175
rect 50725 95147 50759 95175
rect 50787 95147 50821 95175
rect 50849 95147 50883 95175
rect 50911 95147 50959 95175
rect 50649 95113 50959 95147
rect 50649 95085 50697 95113
rect 50725 95085 50759 95113
rect 50787 95085 50821 95113
rect 50849 95085 50883 95113
rect 50911 95085 50959 95113
rect 50649 95051 50959 95085
rect 50649 95023 50697 95051
rect 50725 95023 50759 95051
rect 50787 95023 50821 95051
rect 50849 95023 50883 95051
rect 50911 95023 50959 95051
rect 50649 94989 50959 95023
rect 50649 94961 50697 94989
rect 50725 94961 50759 94989
rect 50787 94961 50821 94989
rect 50849 94961 50883 94989
rect 50911 94961 50959 94989
rect 50649 90103 50959 94961
rect 54624 95175 54784 95192
rect 54624 95147 54659 95175
rect 54687 95147 54721 95175
rect 54749 95147 54784 95175
rect 54624 95113 54784 95147
rect 54624 95085 54659 95113
rect 54687 95085 54721 95113
rect 54749 95085 54784 95113
rect 54624 95051 54784 95085
rect 54624 95023 54659 95051
rect 54687 95023 54721 95051
rect 54749 95023 54784 95051
rect 54624 94989 54784 95023
rect 54624 94961 54659 94989
rect 54687 94961 54721 94989
rect 54749 94961 54784 94989
rect 54624 94944 54784 94961
rect 62304 92175 62464 92192
rect 62304 92147 62339 92175
rect 62367 92147 62401 92175
rect 62429 92147 62464 92175
rect 62304 92113 62464 92147
rect 62304 92085 62339 92113
rect 62367 92085 62401 92113
rect 62429 92085 62464 92113
rect 62304 92051 62464 92085
rect 62304 92023 62339 92051
rect 62367 92023 62401 92051
rect 62429 92023 62464 92051
rect 62304 91989 62464 92023
rect 62304 91961 62339 91989
rect 62367 91961 62401 91989
rect 62429 91961 62464 91989
rect 62304 91944 62464 91961
rect 64149 92175 64459 100961
rect 64149 92147 64197 92175
rect 64225 92147 64259 92175
rect 64287 92147 64321 92175
rect 64349 92147 64383 92175
rect 64411 92147 64459 92175
rect 64149 92113 64459 92147
rect 64149 92085 64197 92113
rect 64225 92085 64259 92113
rect 64287 92085 64321 92113
rect 64349 92085 64383 92113
rect 64411 92085 64459 92113
rect 64149 92051 64459 92085
rect 64149 92023 64197 92051
rect 64225 92023 64259 92051
rect 64287 92023 64321 92051
rect 64349 92023 64383 92051
rect 64411 92023 64459 92051
rect 64149 91989 64459 92023
rect 64149 91961 64197 91989
rect 64225 91961 64259 91989
rect 64287 91961 64321 91989
rect 64349 91961 64383 91989
rect 64411 91961 64459 91989
rect 64149 90103 64459 91961
rect 66009 167175 66319 170745
rect 66009 167147 66057 167175
rect 66085 167147 66119 167175
rect 66147 167147 66181 167175
rect 66209 167147 66243 167175
rect 66271 167147 66319 167175
rect 66009 167113 66319 167147
rect 66009 167085 66057 167113
rect 66085 167085 66119 167113
rect 66147 167085 66181 167113
rect 66209 167085 66243 167113
rect 66271 167085 66319 167113
rect 66009 167051 66319 167085
rect 66009 167023 66057 167051
rect 66085 167023 66119 167051
rect 66147 167023 66181 167051
rect 66209 167023 66243 167051
rect 66271 167023 66319 167051
rect 66009 166989 66319 167023
rect 66009 166961 66057 166989
rect 66085 166961 66119 166989
rect 66147 166961 66181 166989
rect 66209 166961 66243 166989
rect 66271 166961 66319 166989
rect 66009 158175 66319 166961
rect 79509 164175 79819 170745
rect 79509 164147 79557 164175
rect 79585 164147 79619 164175
rect 79647 164147 79681 164175
rect 79709 164147 79743 164175
rect 79771 164147 79819 164175
rect 79509 164113 79819 164147
rect 79509 164085 79557 164113
rect 79585 164085 79619 164113
rect 79647 164085 79681 164113
rect 79709 164085 79743 164113
rect 79771 164085 79819 164113
rect 79509 164051 79819 164085
rect 79509 164023 79557 164051
rect 79585 164023 79619 164051
rect 79647 164023 79681 164051
rect 79709 164023 79743 164051
rect 79771 164023 79819 164051
rect 79509 163989 79819 164023
rect 79509 163961 79557 163989
rect 79585 163961 79619 163989
rect 79647 163961 79681 163989
rect 79709 163961 79743 163989
rect 79771 163961 79819 163989
rect 66009 158147 66057 158175
rect 66085 158147 66119 158175
rect 66147 158147 66181 158175
rect 66209 158147 66243 158175
rect 66271 158147 66319 158175
rect 66009 158113 66319 158147
rect 66009 158085 66057 158113
rect 66085 158085 66119 158113
rect 66147 158085 66181 158113
rect 66209 158085 66243 158113
rect 66271 158085 66319 158113
rect 66009 158051 66319 158085
rect 66009 158023 66057 158051
rect 66085 158023 66119 158051
rect 66147 158023 66181 158051
rect 66209 158023 66243 158051
rect 66271 158023 66319 158051
rect 66009 157989 66319 158023
rect 66009 157961 66057 157989
rect 66085 157961 66119 157989
rect 66147 157961 66181 157989
rect 66209 157961 66243 157989
rect 66271 157961 66319 157989
rect 66009 149175 66319 157961
rect 70624 158175 70784 158192
rect 70624 158147 70659 158175
rect 70687 158147 70721 158175
rect 70749 158147 70784 158175
rect 70624 158113 70784 158147
rect 70624 158085 70659 158113
rect 70687 158085 70721 158113
rect 70749 158085 70784 158113
rect 70624 158051 70784 158085
rect 70624 158023 70659 158051
rect 70687 158023 70721 158051
rect 70749 158023 70784 158051
rect 70624 157989 70784 158023
rect 70624 157961 70659 157989
rect 70687 157961 70721 157989
rect 70749 157961 70784 157989
rect 70624 157944 70784 157961
rect 78304 155175 78464 155192
rect 78304 155147 78339 155175
rect 78367 155147 78401 155175
rect 78429 155147 78464 155175
rect 78304 155113 78464 155147
rect 78304 155085 78339 155113
rect 78367 155085 78401 155113
rect 78429 155085 78464 155113
rect 78304 155051 78464 155085
rect 78304 155023 78339 155051
rect 78367 155023 78401 155051
rect 78429 155023 78464 155051
rect 78304 154989 78464 155023
rect 78304 154961 78339 154989
rect 78367 154961 78401 154989
rect 78429 154961 78464 154989
rect 78304 154944 78464 154961
rect 79509 155175 79819 163961
rect 79509 155147 79557 155175
rect 79585 155147 79619 155175
rect 79647 155147 79681 155175
rect 79709 155147 79743 155175
rect 79771 155147 79819 155175
rect 79509 155113 79819 155147
rect 79509 155085 79557 155113
rect 79585 155085 79619 155113
rect 79647 155085 79681 155113
rect 79709 155085 79743 155113
rect 79771 155085 79819 155113
rect 79509 155051 79819 155085
rect 79509 155023 79557 155051
rect 79585 155023 79619 155051
rect 79647 155023 79681 155051
rect 79709 155023 79743 155051
rect 79771 155023 79819 155051
rect 79509 154989 79819 155023
rect 79509 154961 79557 154989
rect 79585 154961 79619 154989
rect 79647 154961 79681 154989
rect 79709 154961 79743 154989
rect 79771 154961 79819 154989
rect 66009 149147 66057 149175
rect 66085 149147 66119 149175
rect 66147 149147 66181 149175
rect 66209 149147 66243 149175
rect 66271 149147 66319 149175
rect 66009 149113 66319 149147
rect 66009 149085 66057 149113
rect 66085 149085 66119 149113
rect 66147 149085 66181 149113
rect 66209 149085 66243 149113
rect 66271 149085 66319 149113
rect 66009 149051 66319 149085
rect 66009 149023 66057 149051
rect 66085 149023 66119 149051
rect 66147 149023 66181 149051
rect 66209 149023 66243 149051
rect 66271 149023 66319 149051
rect 66009 148989 66319 149023
rect 66009 148961 66057 148989
rect 66085 148961 66119 148989
rect 66147 148961 66181 148989
rect 66209 148961 66243 148989
rect 66271 148961 66319 148989
rect 66009 140175 66319 148961
rect 70624 149175 70784 149192
rect 70624 149147 70659 149175
rect 70687 149147 70721 149175
rect 70749 149147 70784 149175
rect 70624 149113 70784 149147
rect 70624 149085 70659 149113
rect 70687 149085 70721 149113
rect 70749 149085 70784 149113
rect 70624 149051 70784 149085
rect 70624 149023 70659 149051
rect 70687 149023 70721 149051
rect 70749 149023 70784 149051
rect 70624 148989 70784 149023
rect 70624 148961 70659 148989
rect 70687 148961 70721 148989
rect 70749 148961 70784 148989
rect 70624 148944 70784 148961
rect 78304 146175 78464 146192
rect 78304 146147 78339 146175
rect 78367 146147 78401 146175
rect 78429 146147 78464 146175
rect 78304 146113 78464 146147
rect 78304 146085 78339 146113
rect 78367 146085 78401 146113
rect 78429 146085 78464 146113
rect 78304 146051 78464 146085
rect 78304 146023 78339 146051
rect 78367 146023 78401 146051
rect 78429 146023 78464 146051
rect 78304 145989 78464 146023
rect 78304 145961 78339 145989
rect 78367 145961 78401 145989
rect 78429 145961 78464 145989
rect 78304 145944 78464 145961
rect 79509 146175 79819 154961
rect 79509 146147 79557 146175
rect 79585 146147 79619 146175
rect 79647 146147 79681 146175
rect 79709 146147 79743 146175
rect 79771 146147 79819 146175
rect 79509 146113 79819 146147
rect 79509 146085 79557 146113
rect 79585 146085 79619 146113
rect 79647 146085 79681 146113
rect 79709 146085 79743 146113
rect 79771 146085 79819 146113
rect 79509 146051 79819 146085
rect 79509 146023 79557 146051
rect 79585 146023 79619 146051
rect 79647 146023 79681 146051
rect 79709 146023 79743 146051
rect 79771 146023 79819 146051
rect 79509 145989 79819 146023
rect 79509 145961 79557 145989
rect 79585 145961 79619 145989
rect 79647 145961 79681 145989
rect 79709 145961 79743 145989
rect 79771 145961 79819 145989
rect 66009 140147 66057 140175
rect 66085 140147 66119 140175
rect 66147 140147 66181 140175
rect 66209 140147 66243 140175
rect 66271 140147 66319 140175
rect 66009 140113 66319 140147
rect 66009 140085 66057 140113
rect 66085 140085 66119 140113
rect 66147 140085 66181 140113
rect 66209 140085 66243 140113
rect 66271 140085 66319 140113
rect 66009 140051 66319 140085
rect 66009 140023 66057 140051
rect 66085 140023 66119 140051
rect 66147 140023 66181 140051
rect 66209 140023 66243 140051
rect 66271 140023 66319 140051
rect 66009 139989 66319 140023
rect 66009 139961 66057 139989
rect 66085 139961 66119 139989
rect 66147 139961 66181 139989
rect 66209 139961 66243 139989
rect 66271 139961 66319 139989
rect 66009 131175 66319 139961
rect 70624 140175 70784 140192
rect 70624 140147 70659 140175
rect 70687 140147 70721 140175
rect 70749 140147 70784 140175
rect 70624 140113 70784 140147
rect 70624 140085 70659 140113
rect 70687 140085 70721 140113
rect 70749 140085 70784 140113
rect 70624 140051 70784 140085
rect 70624 140023 70659 140051
rect 70687 140023 70721 140051
rect 70749 140023 70784 140051
rect 70624 139989 70784 140023
rect 70624 139961 70659 139989
rect 70687 139961 70721 139989
rect 70749 139961 70784 139989
rect 70624 139944 70784 139961
rect 78304 137175 78464 137192
rect 78304 137147 78339 137175
rect 78367 137147 78401 137175
rect 78429 137147 78464 137175
rect 78304 137113 78464 137147
rect 78304 137085 78339 137113
rect 78367 137085 78401 137113
rect 78429 137085 78464 137113
rect 78304 137051 78464 137085
rect 78304 137023 78339 137051
rect 78367 137023 78401 137051
rect 78429 137023 78464 137051
rect 78304 136989 78464 137023
rect 78304 136961 78339 136989
rect 78367 136961 78401 136989
rect 78429 136961 78464 136989
rect 78304 136944 78464 136961
rect 79509 137175 79819 145961
rect 79509 137147 79557 137175
rect 79585 137147 79619 137175
rect 79647 137147 79681 137175
rect 79709 137147 79743 137175
rect 79771 137147 79819 137175
rect 79509 137113 79819 137147
rect 79509 137085 79557 137113
rect 79585 137085 79619 137113
rect 79647 137085 79681 137113
rect 79709 137085 79743 137113
rect 79771 137085 79819 137113
rect 79509 137051 79819 137085
rect 79509 137023 79557 137051
rect 79585 137023 79619 137051
rect 79647 137023 79681 137051
rect 79709 137023 79743 137051
rect 79771 137023 79819 137051
rect 79509 136989 79819 137023
rect 79509 136961 79557 136989
rect 79585 136961 79619 136989
rect 79647 136961 79681 136989
rect 79709 136961 79743 136989
rect 79771 136961 79819 136989
rect 66009 131147 66057 131175
rect 66085 131147 66119 131175
rect 66147 131147 66181 131175
rect 66209 131147 66243 131175
rect 66271 131147 66319 131175
rect 66009 131113 66319 131147
rect 66009 131085 66057 131113
rect 66085 131085 66119 131113
rect 66147 131085 66181 131113
rect 66209 131085 66243 131113
rect 66271 131085 66319 131113
rect 66009 131051 66319 131085
rect 66009 131023 66057 131051
rect 66085 131023 66119 131051
rect 66147 131023 66181 131051
rect 66209 131023 66243 131051
rect 66271 131023 66319 131051
rect 66009 130989 66319 131023
rect 66009 130961 66057 130989
rect 66085 130961 66119 130989
rect 66147 130961 66181 130989
rect 66209 130961 66243 130989
rect 66271 130961 66319 130989
rect 66009 122175 66319 130961
rect 66009 122147 66057 122175
rect 66085 122147 66119 122175
rect 66147 122147 66181 122175
rect 66209 122147 66243 122175
rect 66271 122147 66319 122175
rect 66009 122113 66319 122147
rect 66009 122085 66057 122113
rect 66085 122085 66119 122113
rect 66147 122085 66181 122113
rect 66209 122085 66243 122113
rect 66271 122085 66319 122113
rect 66009 122051 66319 122085
rect 66009 122023 66057 122051
rect 66085 122023 66119 122051
rect 66147 122023 66181 122051
rect 66209 122023 66243 122051
rect 66271 122023 66319 122051
rect 66009 121989 66319 122023
rect 66009 121961 66057 121989
rect 66085 121961 66119 121989
rect 66147 121961 66181 121989
rect 66209 121961 66243 121989
rect 66271 121961 66319 121989
rect 66009 113175 66319 121961
rect 66009 113147 66057 113175
rect 66085 113147 66119 113175
rect 66147 113147 66181 113175
rect 66209 113147 66243 113175
rect 66271 113147 66319 113175
rect 66009 113113 66319 113147
rect 66009 113085 66057 113113
rect 66085 113085 66119 113113
rect 66147 113085 66181 113113
rect 66209 113085 66243 113113
rect 66271 113085 66319 113113
rect 66009 113051 66319 113085
rect 66009 113023 66057 113051
rect 66085 113023 66119 113051
rect 66147 113023 66181 113051
rect 66209 113023 66243 113051
rect 66271 113023 66319 113051
rect 66009 112989 66319 113023
rect 66009 112961 66057 112989
rect 66085 112961 66119 112989
rect 66147 112961 66181 112989
rect 66209 112961 66243 112989
rect 66271 112961 66319 112989
rect 66009 104175 66319 112961
rect 66009 104147 66057 104175
rect 66085 104147 66119 104175
rect 66147 104147 66181 104175
rect 66209 104147 66243 104175
rect 66271 104147 66319 104175
rect 66009 104113 66319 104147
rect 66009 104085 66057 104113
rect 66085 104085 66119 104113
rect 66147 104085 66181 104113
rect 66209 104085 66243 104113
rect 66271 104085 66319 104113
rect 66009 104051 66319 104085
rect 66009 104023 66057 104051
rect 66085 104023 66119 104051
rect 66147 104023 66181 104051
rect 66209 104023 66243 104051
rect 66271 104023 66319 104051
rect 66009 103989 66319 104023
rect 66009 103961 66057 103989
rect 66085 103961 66119 103989
rect 66147 103961 66181 103989
rect 66209 103961 66243 103989
rect 66271 103961 66319 103989
rect 66009 95175 66319 103961
rect 79509 128175 79819 136961
rect 79509 128147 79557 128175
rect 79585 128147 79619 128175
rect 79647 128147 79681 128175
rect 79709 128147 79743 128175
rect 79771 128147 79819 128175
rect 79509 128113 79819 128147
rect 79509 128085 79557 128113
rect 79585 128085 79619 128113
rect 79647 128085 79681 128113
rect 79709 128085 79743 128113
rect 79771 128085 79819 128113
rect 79509 128051 79819 128085
rect 79509 128023 79557 128051
rect 79585 128023 79619 128051
rect 79647 128023 79681 128051
rect 79709 128023 79743 128051
rect 79771 128023 79819 128051
rect 79509 127989 79819 128023
rect 79509 127961 79557 127989
rect 79585 127961 79619 127989
rect 79647 127961 79681 127989
rect 79709 127961 79743 127989
rect 79771 127961 79819 127989
rect 79509 119175 79819 127961
rect 79509 119147 79557 119175
rect 79585 119147 79619 119175
rect 79647 119147 79681 119175
rect 79709 119147 79743 119175
rect 79771 119147 79819 119175
rect 79509 119113 79819 119147
rect 79509 119085 79557 119113
rect 79585 119085 79619 119113
rect 79647 119085 79681 119113
rect 79709 119085 79743 119113
rect 79771 119085 79819 119113
rect 79509 119051 79819 119085
rect 79509 119023 79557 119051
rect 79585 119023 79619 119051
rect 79647 119023 79681 119051
rect 79709 119023 79743 119051
rect 79771 119023 79819 119051
rect 79509 118989 79819 119023
rect 79509 118961 79557 118989
rect 79585 118961 79619 118989
rect 79647 118961 79681 118989
rect 79709 118961 79743 118989
rect 79771 118961 79819 118989
rect 79509 110175 79819 118961
rect 79509 110147 79557 110175
rect 79585 110147 79619 110175
rect 79647 110147 79681 110175
rect 79709 110147 79743 110175
rect 79771 110147 79819 110175
rect 79509 110113 79819 110147
rect 79509 110085 79557 110113
rect 79585 110085 79619 110113
rect 79647 110085 79681 110113
rect 79709 110085 79743 110113
rect 79771 110085 79819 110113
rect 79509 110051 79819 110085
rect 79509 110023 79557 110051
rect 79585 110023 79619 110051
rect 79647 110023 79681 110051
rect 79709 110023 79743 110051
rect 79771 110023 79819 110051
rect 79509 109989 79819 110023
rect 79509 109961 79557 109989
rect 79585 109961 79619 109989
rect 79647 109961 79681 109989
rect 79709 109961 79743 109989
rect 79771 109961 79819 109989
rect 77664 101175 77824 101192
rect 77664 101147 77699 101175
rect 77727 101147 77761 101175
rect 77789 101147 77824 101175
rect 77664 101113 77824 101147
rect 77664 101085 77699 101113
rect 77727 101085 77761 101113
rect 77789 101085 77824 101113
rect 77664 101051 77824 101085
rect 77664 101023 77699 101051
rect 77727 101023 77761 101051
rect 77789 101023 77824 101051
rect 77664 100989 77824 101023
rect 77664 100961 77699 100989
rect 77727 100961 77761 100989
rect 77789 100961 77824 100989
rect 77664 100944 77824 100961
rect 79509 101175 79819 109961
rect 79509 101147 79557 101175
rect 79585 101147 79619 101175
rect 79647 101147 79681 101175
rect 79709 101147 79743 101175
rect 79771 101147 79819 101175
rect 79509 101113 79819 101147
rect 79509 101085 79557 101113
rect 79585 101085 79619 101113
rect 79647 101085 79681 101113
rect 79709 101085 79743 101113
rect 79771 101085 79819 101113
rect 79509 101051 79819 101085
rect 79509 101023 79557 101051
rect 79585 101023 79619 101051
rect 79647 101023 79681 101051
rect 79709 101023 79743 101051
rect 79771 101023 79819 101051
rect 79509 100989 79819 101023
rect 79509 100961 79557 100989
rect 79585 100961 79619 100989
rect 79647 100961 79681 100989
rect 79709 100961 79743 100989
rect 79771 100961 79819 100989
rect 66009 95147 66057 95175
rect 66085 95147 66119 95175
rect 66147 95147 66181 95175
rect 66209 95147 66243 95175
rect 66271 95147 66319 95175
rect 66009 95113 66319 95147
rect 66009 95085 66057 95113
rect 66085 95085 66119 95113
rect 66147 95085 66181 95113
rect 66209 95085 66243 95113
rect 66271 95085 66319 95113
rect 66009 95051 66319 95085
rect 66009 95023 66057 95051
rect 66085 95023 66119 95051
rect 66147 95023 66181 95051
rect 66209 95023 66243 95051
rect 66271 95023 66319 95051
rect 66009 94989 66319 95023
rect 66009 94961 66057 94989
rect 66085 94961 66119 94989
rect 66147 94961 66181 94989
rect 66209 94961 66243 94989
rect 66271 94961 66319 94989
rect 66009 90103 66319 94961
rect 69984 95175 70144 95192
rect 69984 95147 70019 95175
rect 70047 95147 70081 95175
rect 70109 95147 70144 95175
rect 69984 95113 70144 95147
rect 69984 95085 70019 95113
rect 70047 95085 70081 95113
rect 70109 95085 70144 95113
rect 69984 95051 70144 95085
rect 69984 95023 70019 95051
rect 70047 95023 70081 95051
rect 70109 95023 70144 95051
rect 69984 94989 70144 95023
rect 69984 94961 70019 94989
rect 70047 94961 70081 94989
rect 70109 94961 70144 94989
rect 69984 94944 70144 94961
rect 77664 92175 77824 92192
rect 77664 92147 77699 92175
rect 77727 92147 77761 92175
rect 77789 92147 77824 92175
rect 77664 92113 77824 92147
rect 77664 92085 77699 92113
rect 77727 92085 77761 92113
rect 77789 92085 77824 92113
rect 77664 92051 77824 92085
rect 77664 92023 77699 92051
rect 77727 92023 77761 92051
rect 77789 92023 77824 92051
rect 77664 91989 77824 92023
rect 77664 91961 77699 91989
rect 77727 91961 77761 91989
rect 77789 91961 77824 91989
rect 77664 91944 77824 91961
rect 79509 92175 79819 100961
rect 79509 92147 79557 92175
rect 79585 92147 79619 92175
rect 79647 92147 79681 92175
rect 79709 92147 79743 92175
rect 79771 92147 79819 92175
rect 79509 92113 79819 92147
rect 79509 92085 79557 92113
rect 79585 92085 79619 92113
rect 79647 92085 79681 92113
rect 79709 92085 79743 92113
rect 79771 92085 79819 92113
rect 79509 92051 79819 92085
rect 79509 92023 79557 92051
rect 79585 92023 79619 92051
rect 79647 92023 79681 92051
rect 79709 92023 79743 92051
rect 79771 92023 79819 92051
rect 79509 91989 79819 92023
rect 79509 91961 79557 91989
rect 79585 91961 79619 91989
rect 79647 91961 79681 91989
rect 79709 91961 79743 91989
rect 79771 91961 79819 91989
rect 23904 86175 24064 86192
rect 23904 86147 23939 86175
rect 23967 86147 24001 86175
rect 24029 86147 24064 86175
rect 23904 86113 24064 86147
rect 23904 86085 23939 86113
rect 23967 86085 24001 86113
rect 24029 86085 24064 86113
rect 23904 86051 24064 86085
rect 23904 86023 23939 86051
rect 23967 86023 24001 86051
rect 24029 86023 24064 86051
rect 23904 85989 24064 86023
rect 23904 85961 23939 85989
rect 23967 85961 24001 85989
rect 24029 85961 24064 85989
rect 23904 85944 24064 85961
rect 39264 86175 39424 86192
rect 39264 86147 39299 86175
rect 39327 86147 39361 86175
rect 39389 86147 39424 86175
rect 39264 86113 39424 86147
rect 39264 86085 39299 86113
rect 39327 86085 39361 86113
rect 39389 86085 39424 86113
rect 39264 86051 39424 86085
rect 39264 86023 39299 86051
rect 39327 86023 39361 86051
rect 39389 86023 39424 86051
rect 39264 85989 39424 86023
rect 39264 85961 39299 85989
rect 39327 85961 39361 85989
rect 39389 85961 39424 85989
rect 39264 85944 39424 85961
rect 54624 86175 54784 86192
rect 54624 86147 54659 86175
rect 54687 86147 54721 86175
rect 54749 86147 54784 86175
rect 54624 86113 54784 86147
rect 54624 86085 54659 86113
rect 54687 86085 54721 86113
rect 54749 86085 54784 86113
rect 54624 86051 54784 86085
rect 54624 86023 54659 86051
rect 54687 86023 54721 86051
rect 54749 86023 54784 86051
rect 54624 85989 54784 86023
rect 54624 85961 54659 85989
rect 54687 85961 54721 85989
rect 54749 85961 54784 85989
rect 54624 85944 54784 85961
rect 69984 86175 70144 86192
rect 69984 86147 70019 86175
rect 70047 86147 70081 86175
rect 70109 86147 70144 86175
rect 69984 86113 70144 86147
rect 69984 86085 70019 86113
rect 70047 86085 70081 86113
rect 70109 86085 70144 86113
rect 69984 86051 70144 86085
rect 69984 86023 70019 86051
rect 70047 86023 70081 86051
rect 70109 86023 70144 86051
rect 69984 85989 70144 86023
rect 69984 85961 70019 85989
rect 70047 85961 70081 85989
rect 70109 85961 70144 85989
rect 69984 85944 70144 85961
rect 31584 83175 31744 83192
rect 31584 83147 31619 83175
rect 31647 83147 31681 83175
rect 31709 83147 31744 83175
rect 31584 83113 31744 83147
rect 31584 83085 31619 83113
rect 31647 83085 31681 83113
rect 31709 83085 31744 83113
rect 31584 83051 31744 83085
rect 31584 83023 31619 83051
rect 31647 83023 31681 83051
rect 31709 83023 31744 83051
rect 31584 82989 31744 83023
rect 31584 82961 31619 82989
rect 31647 82961 31681 82989
rect 31709 82961 31744 82989
rect 31584 82944 31744 82961
rect 46944 83175 47104 83192
rect 46944 83147 46979 83175
rect 47007 83147 47041 83175
rect 47069 83147 47104 83175
rect 46944 83113 47104 83147
rect 46944 83085 46979 83113
rect 47007 83085 47041 83113
rect 47069 83085 47104 83113
rect 46944 83051 47104 83085
rect 46944 83023 46979 83051
rect 47007 83023 47041 83051
rect 47069 83023 47104 83051
rect 46944 82989 47104 83023
rect 46944 82961 46979 82989
rect 47007 82961 47041 82989
rect 47069 82961 47104 82989
rect 46944 82944 47104 82961
rect 62304 83175 62464 83192
rect 62304 83147 62339 83175
rect 62367 83147 62401 83175
rect 62429 83147 62464 83175
rect 62304 83113 62464 83147
rect 62304 83085 62339 83113
rect 62367 83085 62401 83113
rect 62429 83085 62464 83113
rect 62304 83051 62464 83085
rect 62304 83023 62339 83051
rect 62367 83023 62401 83051
rect 62429 83023 62464 83051
rect 62304 82989 62464 83023
rect 62304 82961 62339 82989
rect 62367 82961 62401 82989
rect 62429 82961 62464 82989
rect 62304 82944 62464 82961
rect 77664 83175 77824 83192
rect 77664 83147 77699 83175
rect 77727 83147 77761 83175
rect 77789 83147 77824 83175
rect 77664 83113 77824 83147
rect 77664 83085 77699 83113
rect 77727 83085 77761 83113
rect 77789 83085 77824 83113
rect 77664 83051 77824 83085
rect 77664 83023 77699 83051
rect 77727 83023 77761 83051
rect 77789 83023 77824 83051
rect 77664 82989 77824 83023
rect 77664 82961 77699 82989
rect 77727 82961 77761 82989
rect 77789 82961 77824 82989
rect 77664 82944 77824 82961
rect 79509 83175 79819 91961
rect 79509 83147 79557 83175
rect 79585 83147 79619 83175
rect 79647 83147 79681 83175
rect 79709 83147 79743 83175
rect 79771 83147 79819 83175
rect 79509 83113 79819 83147
rect 79509 83085 79557 83113
rect 79585 83085 79619 83113
rect 79647 83085 79681 83113
rect 79709 83085 79743 83113
rect 79771 83085 79819 83113
rect 79509 83051 79819 83085
rect 79509 83023 79557 83051
rect 79585 83023 79619 83051
rect 79647 83023 79681 83051
rect 79709 83023 79743 83051
rect 79771 83023 79819 83051
rect 79509 82989 79819 83023
rect 79509 82961 79557 82989
rect 79585 82961 79619 82989
rect 79647 82961 79681 82989
rect 79709 82961 79743 82989
rect 79771 82961 79819 82989
rect 23904 77175 24064 77192
rect 23904 77147 23939 77175
rect 23967 77147 24001 77175
rect 24029 77147 24064 77175
rect 23904 77113 24064 77147
rect 23904 77085 23939 77113
rect 23967 77085 24001 77113
rect 24029 77085 24064 77113
rect 23904 77051 24064 77085
rect 23904 77023 23939 77051
rect 23967 77023 24001 77051
rect 24029 77023 24064 77051
rect 23904 76989 24064 77023
rect 23904 76961 23939 76989
rect 23967 76961 24001 76989
rect 24029 76961 24064 76989
rect 23904 76944 24064 76961
rect 39264 77175 39424 77192
rect 39264 77147 39299 77175
rect 39327 77147 39361 77175
rect 39389 77147 39424 77175
rect 39264 77113 39424 77147
rect 39264 77085 39299 77113
rect 39327 77085 39361 77113
rect 39389 77085 39424 77113
rect 39264 77051 39424 77085
rect 39264 77023 39299 77051
rect 39327 77023 39361 77051
rect 39389 77023 39424 77051
rect 39264 76989 39424 77023
rect 39264 76961 39299 76989
rect 39327 76961 39361 76989
rect 39389 76961 39424 76989
rect 39264 76944 39424 76961
rect 54624 77175 54784 77192
rect 54624 77147 54659 77175
rect 54687 77147 54721 77175
rect 54749 77147 54784 77175
rect 54624 77113 54784 77147
rect 54624 77085 54659 77113
rect 54687 77085 54721 77113
rect 54749 77085 54784 77113
rect 54624 77051 54784 77085
rect 54624 77023 54659 77051
rect 54687 77023 54721 77051
rect 54749 77023 54784 77051
rect 54624 76989 54784 77023
rect 54624 76961 54659 76989
rect 54687 76961 54721 76989
rect 54749 76961 54784 76989
rect 54624 76944 54784 76961
rect 69984 77175 70144 77192
rect 69984 77147 70019 77175
rect 70047 77147 70081 77175
rect 70109 77147 70144 77175
rect 69984 77113 70144 77147
rect 69984 77085 70019 77113
rect 70047 77085 70081 77113
rect 70109 77085 70144 77113
rect 69984 77051 70144 77085
rect 69984 77023 70019 77051
rect 70047 77023 70081 77051
rect 70109 77023 70144 77051
rect 69984 76989 70144 77023
rect 69984 76961 70019 76989
rect 70047 76961 70081 76989
rect 70109 76961 70144 76989
rect 69984 76944 70144 76961
rect 21406 74713 21434 74718
rect 19929 68147 19977 68175
rect 20005 68147 20039 68175
rect 20067 68147 20101 68175
rect 20129 68147 20163 68175
rect 20191 68147 20239 68175
rect 19929 68113 20239 68147
rect 19929 68085 19977 68113
rect 20005 68085 20039 68113
rect 20067 68085 20101 68113
rect 20129 68085 20163 68113
rect 20191 68085 20239 68113
rect 19929 68051 20239 68085
rect 19929 68023 19977 68051
rect 20005 68023 20039 68051
rect 20067 68023 20101 68051
rect 20129 68023 20163 68051
rect 20191 68023 20239 68051
rect 19929 67989 20239 68023
rect 19929 67961 19977 67989
rect 20005 67961 20039 67989
rect 20067 67961 20101 67989
rect 20129 67961 20163 67989
rect 20191 67961 20239 67989
rect 19929 59175 20239 67961
rect 19929 59147 19977 59175
rect 20005 59147 20039 59175
rect 20067 59147 20101 59175
rect 20129 59147 20163 59175
rect 20191 59147 20239 59175
rect 19929 59113 20239 59147
rect 19929 59085 19977 59113
rect 20005 59085 20039 59113
rect 20067 59085 20101 59113
rect 20129 59085 20163 59113
rect 20191 59085 20239 59113
rect 19929 59051 20239 59085
rect 19929 59023 19977 59051
rect 20005 59023 20039 59051
rect 20067 59023 20101 59051
rect 20129 59023 20163 59051
rect 20191 59023 20239 59051
rect 19929 58989 20239 59023
rect 19929 58961 19977 58989
rect 20005 58961 20039 58989
rect 20067 58961 20101 58989
rect 20129 58961 20163 58989
rect 20191 58961 20239 58989
rect 19929 50175 20239 58961
rect 19929 50147 19977 50175
rect 20005 50147 20039 50175
rect 20067 50147 20101 50175
rect 20129 50147 20163 50175
rect 20191 50147 20239 50175
rect 19929 50113 20239 50147
rect 19929 50085 19977 50113
rect 20005 50085 20039 50113
rect 20067 50085 20101 50113
rect 20129 50085 20163 50113
rect 20191 50085 20239 50113
rect 19929 50051 20239 50085
rect 19929 50023 19977 50051
rect 20005 50023 20039 50051
rect 20067 50023 20101 50051
rect 20129 50023 20163 50051
rect 20191 50023 20239 50051
rect 19929 49989 20239 50023
rect 19929 49961 19977 49989
rect 20005 49961 20039 49989
rect 20067 49961 20101 49989
rect 20129 49961 20163 49989
rect 20191 49961 20239 49989
rect 19929 41175 20239 49961
rect 19929 41147 19977 41175
rect 20005 41147 20039 41175
rect 20067 41147 20101 41175
rect 20129 41147 20163 41175
rect 20191 41147 20239 41175
rect 19929 41113 20239 41147
rect 19929 41085 19977 41113
rect 20005 41085 20039 41113
rect 20067 41085 20101 41113
rect 20129 41085 20163 41113
rect 20191 41085 20239 41113
rect 19929 41051 20239 41085
rect 19929 41023 19977 41051
rect 20005 41023 20039 41051
rect 20067 41023 20101 41051
rect 20129 41023 20163 41051
rect 20191 41023 20239 41051
rect 19929 40989 20239 41023
rect 19929 40961 19977 40989
rect 20005 40961 20039 40989
rect 20067 40961 20101 40989
rect 20129 40961 20163 40989
rect 20191 40961 20239 40989
rect 19929 32175 20239 40961
rect 19929 32147 19977 32175
rect 20005 32147 20039 32175
rect 20067 32147 20101 32175
rect 20129 32147 20163 32175
rect 20191 32147 20239 32175
rect 19929 32113 20239 32147
rect 19929 32085 19977 32113
rect 20005 32085 20039 32113
rect 20067 32085 20101 32113
rect 20129 32085 20163 32113
rect 20191 32085 20239 32113
rect 19929 32051 20239 32085
rect 19929 32023 19977 32051
rect 20005 32023 20039 32051
rect 20067 32023 20101 32051
rect 20129 32023 20163 32051
rect 20191 32023 20239 32051
rect 19929 31989 20239 32023
rect 19929 31961 19977 31989
rect 20005 31961 20039 31989
rect 20067 31961 20101 31989
rect 20129 31961 20163 31989
rect 20191 31961 20239 31989
rect 19929 23175 20239 31961
rect 19929 23147 19977 23175
rect 20005 23147 20039 23175
rect 20067 23147 20101 23175
rect 20129 23147 20163 23175
rect 20191 23147 20239 23175
rect 19929 23113 20239 23147
rect 19929 23085 19977 23113
rect 20005 23085 20039 23113
rect 20067 23085 20101 23113
rect 20129 23085 20163 23113
rect 20191 23085 20239 23113
rect 19929 23051 20239 23085
rect 19929 23023 19977 23051
rect 20005 23023 20039 23051
rect 20067 23023 20101 23051
rect 20129 23023 20163 23051
rect 20191 23023 20239 23051
rect 19929 22989 20239 23023
rect 19929 22961 19977 22989
rect 20005 22961 20039 22989
rect 20067 22961 20101 22989
rect 20129 22961 20163 22989
rect 20191 22961 20239 22989
rect 19929 14175 20239 22961
rect 19929 14147 19977 14175
rect 20005 14147 20039 14175
rect 20067 14147 20101 14175
rect 20129 14147 20163 14175
rect 20191 14147 20239 14175
rect 19929 14113 20239 14147
rect 19929 14085 19977 14113
rect 20005 14085 20039 14113
rect 20067 14085 20101 14113
rect 20129 14085 20163 14113
rect 20191 14085 20239 14113
rect 19929 14051 20239 14085
rect 19929 14023 19977 14051
rect 20005 14023 20039 14051
rect 20067 14023 20101 14051
rect 20129 14023 20163 14051
rect 20191 14023 20239 14051
rect 19929 13989 20239 14023
rect 19929 13961 19977 13989
rect 20005 13961 20039 13989
rect 20067 13961 20101 13989
rect 20129 13961 20163 13989
rect 20191 13961 20239 13989
rect 19929 5175 20239 13961
rect 19929 5147 19977 5175
rect 20005 5147 20039 5175
rect 20067 5147 20101 5175
rect 20129 5147 20163 5175
rect 20191 5147 20239 5175
rect 19929 5113 20239 5147
rect 19929 5085 19977 5113
rect 20005 5085 20039 5113
rect 20067 5085 20101 5113
rect 20129 5085 20163 5113
rect 20191 5085 20239 5113
rect 19929 5051 20239 5085
rect 19929 5023 19977 5051
rect 20005 5023 20039 5051
rect 20067 5023 20101 5051
rect 20129 5023 20163 5051
rect 20191 5023 20239 5051
rect 19929 4989 20239 5023
rect 19929 4961 19977 4989
rect 20005 4961 20039 4989
rect 20067 4961 20101 4989
rect 20129 4961 20163 4989
rect 20191 4961 20239 4989
rect 19929 -560 20239 4961
rect 19929 -588 19977 -560
rect 20005 -588 20039 -560
rect 20067 -588 20101 -560
rect 20129 -588 20163 -560
rect 20191 -588 20239 -560
rect 19929 -622 20239 -588
rect 19929 -650 19977 -622
rect 20005 -650 20039 -622
rect 20067 -650 20101 -622
rect 20129 -650 20163 -622
rect 20191 -650 20239 -622
rect 19929 -684 20239 -650
rect 19929 -712 19977 -684
rect 20005 -712 20039 -684
rect 20067 -712 20101 -684
rect 20129 -712 20163 -684
rect 20191 -712 20239 -684
rect 19929 -746 20239 -712
rect 19929 -774 19977 -746
rect 20005 -774 20039 -746
rect 20067 -774 20101 -746
rect 20129 -774 20163 -746
rect 20191 -774 20239 -746
rect 19929 -822 20239 -774
rect 33429 74175 33739 74345
rect 33429 74147 33477 74175
rect 33505 74147 33539 74175
rect 33567 74147 33601 74175
rect 33629 74147 33663 74175
rect 33691 74147 33739 74175
rect 33429 74113 33739 74147
rect 33429 74085 33477 74113
rect 33505 74085 33539 74113
rect 33567 74085 33601 74113
rect 33629 74085 33663 74113
rect 33691 74085 33739 74113
rect 33429 74051 33739 74085
rect 33429 74023 33477 74051
rect 33505 74023 33539 74051
rect 33567 74023 33601 74051
rect 33629 74023 33663 74051
rect 33691 74023 33739 74051
rect 33429 73989 33739 74023
rect 33429 73961 33477 73989
rect 33505 73961 33539 73989
rect 33567 73961 33601 73989
rect 33629 73961 33663 73989
rect 33691 73961 33739 73989
rect 33429 65175 33739 73961
rect 33429 65147 33477 65175
rect 33505 65147 33539 65175
rect 33567 65147 33601 65175
rect 33629 65147 33663 65175
rect 33691 65147 33739 65175
rect 33429 65113 33739 65147
rect 33429 65085 33477 65113
rect 33505 65085 33539 65113
rect 33567 65085 33601 65113
rect 33629 65085 33663 65113
rect 33691 65085 33739 65113
rect 33429 65051 33739 65085
rect 33429 65023 33477 65051
rect 33505 65023 33539 65051
rect 33567 65023 33601 65051
rect 33629 65023 33663 65051
rect 33691 65023 33739 65051
rect 33429 64989 33739 65023
rect 33429 64961 33477 64989
rect 33505 64961 33539 64989
rect 33567 64961 33601 64989
rect 33629 64961 33663 64989
rect 33691 64961 33739 64989
rect 33429 56175 33739 64961
rect 33429 56147 33477 56175
rect 33505 56147 33539 56175
rect 33567 56147 33601 56175
rect 33629 56147 33663 56175
rect 33691 56147 33739 56175
rect 33429 56113 33739 56147
rect 33429 56085 33477 56113
rect 33505 56085 33539 56113
rect 33567 56085 33601 56113
rect 33629 56085 33663 56113
rect 33691 56085 33739 56113
rect 33429 56051 33739 56085
rect 33429 56023 33477 56051
rect 33505 56023 33539 56051
rect 33567 56023 33601 56051
rect 33629 56023 33663 56051
rect 33691 56023 33739 56051
rect 33429 55989 33739 56023
rect 33429 55961 33477 55989
rect 33505 55961 33539 55989
rect 33567 55961 33601 55989
rect 33629 55961 33663 55989
rect 33691 55961 33739 55989
rect 33429 47175 33739 55961
rect 33429 47147 33477 47175
rect 33505 47147 33539 47175
rect 33567 47147 33601 47175
rect 33629 47147 33663 47175
rect 33691 47147 33739 47175
rect 33429 47113 33739 47147
rect 33429 47085 33477 47113
rect 33505 47085 33539 47113
rect 33567 47085 33601 47113
rect 33629 47085 33663 47113
rect 33691 47085 33739 47113
rect 33429 47051 33739 47085
rect 33429 47023 33477 47051
rect 33505 47023 33539 47051
rect 33567 47023 33601 47051
rect 33629 47023 33663 47051
rect 33691 47023 33739 47051
rect 33429 46989 33739 47023
rect 33429 46961 33477 46989
rect 33505 46961 33539 46989
rect 33567 46961 33601 46989
rect 33629 46961 33663 46989
rect 33691 46961 33739 46989
rect 33429 38175 33739 46961
rect 33429 38147 33477 38175
rect 33505 38147 33539 38175
rect 33567 38147 33601 38175
rect 33629 38147 33663 38175
rect 33691 38147 33739 38175
rect 33429 38113 33739 38147
rect 33429 38085 33477 38113
rect 33505 38085 33539 38113
rect 33567 38085 33601 38113
rect 33629 38085 33663 38113
rect 33691 38085 33739 38113
rect 33429 38051 33739 38085
rect 33429 38023 33477 38051
rect 33505 38023 33539 38051
rect 33567 38023 33601 38051
rect 33629 38023 33663 38051
rect 33691 38023 33739 38051
rect 33429 37989 33739 38023
rect 33429 37961 33477 37989
rect 33505 37961 33539 37989
rect 33567 37961 33601 37989
rect 33629 37961 33663 37989
rect 33691 37961 33739 37989
rect 33429 29175 33739 37961
rect 33429 29147 33477 29175
rect 33505 29147 33539 29175
rect 33567 29147 33601 29175
rect 33629 29147 33663 29175
rect 33691 29147 33739 29175
rect 33429 29113 33739 29147
rect 33429 29085 33477 29113
rect 33505 29085 33539 29113
rect 33567 29085 33601 29113
rect 33629 29085 33663 29113
rect 33691 29085 33739 29113
rect 33429 29051 33739 29085
rect 33429 29023 33477 29051
rect 33505 29023 33539 29051
rect 33567 29023 33601 29051
rect 33629 29023 33663 29051
rect 33691 29023 33739 29051
rect 33429 28989 33739 29023
rect 33429 28961 33477 28989
rect 33505 28961 33539 28989
rect 33567 28961 33601 28989
rect 33629 28961 33663 28989
rect 33691 28961 33739 28989
rect 33429 20175 33739 28961
rect 33429 20147 33477 20175
rect 33505 20147 33539 20175
rect 33567 20147 33601 20175
rect 33629 20147 33663 20175
rect 33691 20147 33739 20175
rect 33429 20113 33739 20147
rect 33429 20085 33477 20113
rect 33505 20085 33539 20113
rect 33567 20085 33601 20113
rect 33629 20085 33663 20113
rect 33691 20085 33739 20113
rect 33429 20051 33739 20085
rect 33429 20023 33477 20051
rect 33505 20023 33539 20051
rect 33567 20023 33601 20051
rect 33629 20023 33663 20051
rect 33691 20023 33739 20051
rect 33429 19989 33739 20023
rect 33429 19961 33477 19989
rect 33505 19961 33539 19989
rect 33567 19961 33601 19989
rect 33629 19961 33663 19989
rect 33691 19961 33739 19989
rect 33429 11175 33739 19961
rect 33429 11147 33477 11175
rect 33505 11147 33539 11175
rect 33567 11147 33601 11175
rect 33629 11147 33663 11175
rect 33691 11147 33739 11175
rect 33429 11113 33739 11147
rect 33429 11085 33477 11113
rect 33505 11085 33539 11113
rect 33567 11085 33601 11113
rect 33629 11085 33663 11113
rect 33691 11085 33739 11113
rect 33429 11051 33739 11085
rect 33429 11023 33477 11051
rect 33505 11023 33539 11051
rect 33567 11023 33601 11051
rect 33629 11023 33663 11051
rect 33691 11023 33739 11051
rect 33429 10989 33739 11023
rect 33429 10961 33477 10989
rect 33505 10961 33539 10989
rect 33567 10961 33601 10989
rect 33629 10961 33663 10989
rect 33691 10961 33739 10989
rect 33429 2175 33739 10961
rect 33429 2147 33477 2175
rect 33505 2147 33539 2175
rect 33567 2147 33601 2175
rect 33629 2147 33663 2175
rect 33691 2147 33739 2175
rect 33429 2113 33739 2147
rect 33429 2085 33477 2113
rect 33505 2085 33539 2113
rect 33567 2085 33601 2113
rect 33629 2085 33663 2113
rect 33691 2085 33739 2113
rect 33429 2051 33739 2085
rect 33429 2023 33477 2051
rect 33505 2023 33539 2051
rect 33567 2023 33601 2051
rect 33629 2023 33663 2051
rect 33691 2023 33739 2051
rect 33429 1989 33739 2023
rect 33429 1961 33477 1989
rect 33505 1961 33539 1989
rect 33567 1961 33601 1989
rect 33629 1961 33663 1989
rect 33691 1961 33739 1989
rect 33429 -80 33739 1961
rect 33429 -108 33477 -80
rect 33505 -108 33539 -80
rect 33567 -108 33601 -80
rect 33629 -108 33663 -80
rect 33691 -108 33739 -80
rect 33429 -142 33739 -108
rect 33429 -170 33477 -142
rect 33505 -170 33539 -142
rect 33567 -170 33601 -142
rect 33629 -170 33663 -142
rect 33691 -170 33739 -142
rect 33429 -204 33739 -170
rect 33429 -232 33477 -204
rect 33505 -232 33539 -204
rect 33567 -232 33601 -204
rect 33629 -232 33663 -204
rect 33691 -232 33739 -204
rect 33429 -266 33739 -232
rect 33429 -294 33477 -266
rect 33505 -294 33539 -266
rect 33567 -294 33601 -266
rect 33629 -294 33663 -266
rect 33691 -294 33739 -266
rect 33429 -822 33739 -294
rect 35289 68175 35599 74345
rect 35289 68147 35337 68175
rect 35365 68147 35399 68175
rect 35427 68147 35461 68175
rect 35489 68147 35523 68175
rect 35551 68147 35599 68175
rect 35289 68113 35599 68147
rect 35289 68085 35337 68113
rect 35365 68085 35399 68113
rect 35427 68085 35461 68113
rect 35489 68085 35523 68113
rect 35551 68085 35599 68113
rect 35289 68051 35599 68085
rect 35289 68023 35337 68051
rect 35365 68023 35399 68051
rect 35427 68023 35461 68051
rect 35489 68023 35523 68051
rect 35551 68023 35599 68051
rect 35289 67989 35599 68023
rect 35289 67961 35337 67989
rect 35365 67961 35399 67989
rect 35427 67961 35461 67989
rect 35489 67961 35523 67989
rect 35551 67961 35599 67989
rect 35289 59175 35599 67961
rect 35289 59147 35337 59175
rect 35365 59147 35399 59175
rect 35427 59147 35461 59175
rect 35489 59147 35523 59175
rect 35551 59147 35599 59175
rect 35289 59113 35599 59147
rect 35289 59085 35337 59113
rect 35365 59085 35399 59113
rect 35427 59085 35461 59113
rect 35489 59085 35523 59113
rect 35551 59085 35599 59113
rect 35289 59051 35599 59085
rect 35289 59023 35337 59051
rect 35365 59023 35399 59051
rect 35427 59023 35461 59051
rect 35489 59023 35523 59051
rect 35551 59023 35599 59051
rect 35289 58989 35599 59023
rect 35289 58961 35337 58989
rect 35365 58961 35399 58989
rect 35427 58961 35461 58989
rect 35489 58961 35523 58989
rect 35551 58961 35599 58989
rect 35289 50175 35599 58961
rect 35289 50147 35337 50175
rect 35365 50147 35399 50175
rect 35427 50147 35461 50175
rect 35489 50147 35523 50175
rect 35551 50147 35599 50175
rect 35289 50113 35599 50147
rect 35289 50085 35337 50113
rect 35365 50085 35399 50113
rect 35427 50085 35461 50113
rect 35489 50085 35523 50113
rect 35551 50085 35599 50113
rect 35289 50051 35599 50085
rect 35289 50023 35337 50051
rect 35365 50023 35399 50051
rect 35427 50023 35461 50051
rect 35489 50023 35523 50051
rect 35551 50023 35599 50051
rect 35289 49989 35599 50023
rect 35289 49961 35337 49989
rect 35365 49961 35399 49989
rect 35427 49961 35461 49989
rect 35489 49961 35523 49989
rect 35551 49961 35599 49989
rect 35289 41175 35599 49961
rect 35289 41147 35337 41175
rect 35365 41147 35399 41175
rect 35427 41147 35461 41175
rect 35489 41147 35523 41175
rect 35551 41147 35599 41175
rect 35289 41113 35599 41147
rect 35289 41085 35337 41113
rect 35365 41085 35399 41113
rect 35427 41085 35461 41113
rect 35489 41085 35523 41113
rect 35551 41085 35599 41113
rect 35289 41051 35599 41085
rect 35289 41023 35337 41051
rect 35365 41023 35399 41051
rect 35427 41023 35461 41051
rect 35489 41023 35523 41051
rect 35551 41023 35599 41051
rect 35289 40989 35599 41023
rect 35289 40961 35337 40989
rect 35365 40961 35399 40989
rect 35427 40961 35461 40989
rect 35489 40961 35523 40989
rect 35551 40961 35599 40989
rect 35289 32175 35599 40961
rect 35289 32147 35337 32175
rect 35365 32147 35399 32175
rect 35427 32147 35461 32175
rect 35489 32147 35523 32175
rect 35551 32147 35599 32175
rect 35289 32113 35599 32147
rect 35289 32085 35337 32113
rect 35365 32085 35399 32113
rect 35427 32085 35461 32113
rect 35489 32085 35523 32113
rect 35551 32085 35599 32113
rect 35289 32051 35599 32085
rect 35289 32023 35337 32051
rect 35365 32023 35399 32051
rect 35427 32023 35461 32051
rect 35489 32023 35523 32051
rect 35551 32023 35599 32051
rect 35289 31989 35599 32023
rect 35289 31961 35337 31989
rect 35365 31961 35399 31989
rect 35427 31961 35461 31989
rect 35489 31961 35523 31989
rect 35551 31961 35599 31989
rect 35289 23175 35599 31961
rect 35289 23147 35337 23175
rect 35365 23147 35399 23175
rect 35427 23147 35461 23175
rect 35489 23147 35523 23175
rect 35551 23147 35599 23175
rect 35289 23113 35599 23147
rect 35289 23085 35337 23113
rect 35365 23085 35399 23113
rect 35427 23085 35461 23113
rect 35489 23085 35523 23113
rect 35551 23085 35599 23113
rect 35289 23051 35599 23085
rect 35289 23023 35337 23051
rect 35365 23023 35399 23051
rect 35427 23023 35461 23051
rect 35489 23023 35523 23051
rect 35551 23023 35599 23051
rect 35289 22989 35599 23023
rect 35289 22961 35337 22989
rect 35365 22961 35399 22989
rect 35427 22961 35461 22989
rect 35489 22961 35523 22989
rect 35551 22961 35599 22989
rect 35289 14175 35599 22961
rect 35289 14147 35337 14175
rect 35365 14147 35399 14175
rect 35427 14147 35461 14175
rect 35489 14147 35523 14175
rect 35551 14147 35599 14175
rect 35289 14113 35599 14147
rect 35289 14085 35337 14113
rect 35365 14085 35399 14113
rect 35427 14085 35461 14113
rect 35489 14085 35523 14113
rect 35551 14085 35599 14113
rect 35289 14051 35599 14085
rect 35289 14023 35337 14051
rect 35365 14023 35399 14051
rect 35427 14023 35461 14051
rect 35489 14023 35523 14051
rect 35551 14023 35599 14051
rect 35289 13989 35599 14023
rect 35289 13961 35337 13989
rect 35365 13961 35399 13989
rect 35427 13961 35461 13989
rect 35489 13961 35523 13989
rect 35551 13961 35599 13989
rect 35289 5175 35599 13961
rect 35289 5147 35337 5175
rect 35365 5147 35399 5175
rect 35427 5147 35461 5175
rect 35489 5147 35523 5175
rect 35551 5147 35599 5175
rect 35289 5113 35599 5147
rect 35289 5085 35337 5113
rect 35365 5085 35399 5113
rect 35427 5085 35461 5113
rect 35489 5085 35523 5113
rect 35551 5085 35599 5113
rect 35289 5051 35599 5085
rect 35289 5023 35337 5051
rect 35365 5023 35399 5051
rect 35427 5023 35461 5051
rect 35489 5023 35523 5051
rect 35551 5023 35599 5051
rect 35289 4989 35599 5023
rect 35289 4961 35337 4989
rect 35365 4961 35399 4989
rect 35427 4961 35461 4989
rect 35489 4961 35523 4989
rect 35551 4961 35599 4989
rect 35289 -560 35599 4961
rect 35289 -588 35337 -560
rect 35365 -588 35399 -560
rect 35427 -588 35461 -560
rect 35489 -588 35523 -560
rect 35551 -588 35599 -560
rect 35289 -622 35599 -588
rect 35289 -650 35337 -622
rect 35365 -650 35399 -622
rect 35427 -650 35461 -622
rect 35489 -650 35523 -622
rect 35551 -650 35599 -622
rect 35289 -684 35599 -650
rect 35289 -712 35337 -684
rect 35365 -712 35399 -684
rect 35427 -712 35461 -684
rect 35489 -712 35523 -684
rect 35551 -712 35599 -684
rect 35289 -746 35599 -712
rect 35289 -774 35337 -746
rect 35365 -774 35399 -746
rect 35427 -774 35461 -746
rect 35489 -774 35523 -746
rect 35551 -774 35599 -746
rect 35289 -822 35599 -774
rect 48789 74175 49099 74345
rect 48789 74147 48837 74175
rect 48865 74147 48899 74175
rect 48927 74147 48961 74175
rect 48989 74147 49023 74175
rect 49051 74147 49099 74175
rect 48789 74113 49099 74147
rect 48789 74085 48837 74113
rect 48865 74085 48899 74113
rect 48927 74085 48961 74113
rect 48989 74085 49023 74113
rect 49051 74085 49099 74113
rect 48789 74051 49099 74085
rect 48789 74023 48837 74051
rect 48865 74023 48899 74051
rect 48927 74023 48961 74051
rect 48989 74023 49023 74051
rect 49051 74023 49099 74051
rect 48789 73989 49099 74023
rect 48789 73961 48837 73989
rect 48865 73961 48899 73989
rect 48927 73961 48961 73989
rect 48989 73961 49023 73989
rect 49051 73961 49099 73989
rect 48789 65175 49099 73961
rect 48789 65147 48837 65175
rect 48865 65147 48899 65175
rect 48927 65147 48961 65175
rect 48989 65147 49023 65175
rect 49051 65147 49099 65175
rect 48789 65113 49099 65147
rect 48789 65085 48837 65113
rect 48865 65085 48899 65113
rect 48927 65085 48961 65113
rect 48989 65085 49023 65113
rect 49051 65085 49099 65113
rect 48789 65051 49099 65085
rect 48789 65023 48837 65051
rect 48865 65023 48899 65051
rect 48927 65023 48961 65051
rect 48989 65023 49023 65051
rect 49051 65023 49099 65051
rect 48789 64989 49099 65023
rect 48789 64961 48837 64989
rect 48865 64961 48899 64989
rect 48927 64961 48961 64989
rect 48989 64961 49023 64989
rect 49051 64961 49099 64989
rect 48789 56175 49099 64961
rect 48789 56147 48837 56175
rect 48865 56147 48899 56175
rect 48927 56147 48961 56175
rect 48989 56147 49023 56175
rect 49051 56147 49099 56175
rect 48789 56113 49099 56147
rect 48789 56085 48837 56113
rect 48865 56085 48899 56113
rect 48927 56085 48961 56113
rect 48989 56085 49023 56113
rect 49051 56085 49099 56113
rect 48789 56051 49099 56085
rect 48789 56023 48837 56051
rect 48865 56023 48899 56051
rect 48927 56023 48961 56051
rect 48989 56023 49023 56051
rect 49051 56023 49099 56051
rect 48789 55989 49099 56023
rect 48789 55961 48837 55989
rect 48865 55961 48899 55989
rect 48927 55961 48961 55989
rect 48989 55961 49023 55989
rect 49051 55961 49099 55989
rect 48789 47175 49099 55961
rect 48789 47147 48837 47175
rect 48865 47147 48899 47175
rect 48927 47147 48961 47175
rect 48989 47147 49023 47175
rect 49051 47147 49099 47175
rect 48789 47113 49099 47147
rect 48789 47085 48837 47113
rect 48865 47085 48899 47113
rect 48927 47085 48961 47113
rect 48989 47085 49023 47113
rect 49051 47085 49099 47113
rect 48789 47051 49099 47085
rect 48789 47023 48837 47051
rect 48865 47023 48899 47051
rect 48927 47023 48961 47051
rect 48989 47023 49023 47051
rect 49051 47023 49099 47051
rect 48789 46989 49099 47023
rect 48789 46961 48837 46989
rect 48865 46961 48899 46989
rect 48927 46961 48961 46989
rect 48989 46961 49023 46989
rect 49051 46961 49099 46989
rect 48789 38175 49099 46961
rect 48789 38147 48837 38175
rect 48865 38147 48899 38175
rect 48927 38147 48961 38175
rect 48989 38147 49023 38175
rect 49051 38147 49099 38175
rect 48789 38113 49099 38147
rect 48789 38085 48837 38113
rect 48865 38085 48899 38113
rect 48927 38085 48961 38113
rect 48989 38085 49023 38113
rect 49051 38085 49099 38113
rect 48789 38051 49099 38085
rect 48789 38023 48837 38051
rect 48865 38023 48899 38051
rect 48927 38023 48961 38051
rect 48989 38023 49023 38051
rect 49051 38023 49099 38051
rect 48789 37989 49099 38023
rect 48789 37961 48837 37989
rect 48865 37961 48899 37989
rect 48927 37961 48961 37989
rect 48989 37961 49023 37989
rect 49051 37961 49099 37989
rect 48789 29175 49099 37961
rect 48789 29147 48837 29175
rect 48865 29147 48899 29175
rect 48927 29147 48961 29175
rect 48989 29147 49023 29175
rect 49051 29147 49099 29175
rect 48789 29113 49099 29147
rect 48789 29085 48837 29113
rect 48865 29085 48899 29113
rect 48927 29085 48961 29113
rect 48989 29085 49023 29113
rect 49051 29085 49099 29113
rect 48789 29051 49099 29085
rect 48789 29023 48837 29051
rect 48865 29023 48899 29051
rect 48927 29023 48961 29051
rect 48989 29023 49023 29051
rect 49051 29023 49099 29051
rect 48789 28989 49099 29023
rect 48789 28961 48837 28989
rect 48865 28961 48899 28989
rect 48927 28961 48961 28989
rect 48989 28961 49023 28989
rect 49051 28961 49099 28989
rect 48789 20175 49099 28961
rect 48789 20147 48837 20175
rect 48865 20147 48899 20175
rect 48927 20147 48961 20175
rect 48989 20147 49023 20175
rect 49051 20147 49099 20175
rect 48789 20113 49099 20147
rect 48789 20085 48837 20113
rect 48865 20085 48899 20113
rect 48927 20085 48961 20113
rect 48989 20085 49023 20113
rect 49051 20085 49099 20113
rect 48789 20051 49099 20085
rect 48789 20023 48837 20051
rect 48865 20023 48899 20051
rect 48927 20023 48961 20051
rect 48989 20023 49023 20051
rect 49051 20023 49099 20051
rect 48789 19989 49099 20023
rect 48789 19961 48837 19989
rect 48865 19961 48899 19989
rect 48927 19961 48961 19989
rect 48989 19961 49023 19989
rect 49051 19961 49099 19989
rect 48789 11175 49099 19961
rect 48789 11147 48837 11175
rect 48865 11147 48899 11175
rect 48927 11147 48961 11175
rect 48989 11147 49023 11175
rect 49051 11147 49099 11175
rect 48789 11113 49099 11147
rect 48789 11085 48837 11113
rect 48865 11085 48899 11113
rect 48927 11085 48961 11113
rect 48989 11085 49023 11113
rect 49051 11085 49099 11113
rect 48789 11051 49099 11085
rect 48789 11023 48837 11051
rect 48865 11023 48899 11051
rect 48927 11023 48961 11051
rect 48989 11023 49023 11051
rect 49051 11023 49099 11051
rect 48789 10989 49099 11023
rect 48789 10961 48837 10989
rect 48865 10961 48899 10989
rect 48927 10961 48961 10989
rect 48989 10961 49023 10989
rect 49051 10961 49099 10989
rect 48789 2175 49099 10961
rect 48789 2147 48837 2175
rect 48865 2147 48899 2175
rect 48927 2147 48961 2175
rect 48989 2147 49023 2175
rect 49051 2147 49099 2175
rect 48789 2113 49099 2147
rect 48789 2085 48837 2113
rect 48865 2085 48899 2113
rect 48927 2085 48961 2113
rect 48989 2085 49023 2113
rect 49051 2085 49099 2113
rect 48789 2051 49099 2085
rect 48789 2023 48837 2051
rect 48865 2023 48899 2051
rect 48927 2023 48961 2051
rect 48989 2023 49023 2051
rect 49051 2023 49099 2051
rect 48789 1989 49099 2023
rect 48789 1961 48837 1989
rect 48865 1961 48899 1989
rect 48927 1961 48961 1989
rect 48989 1961 49023 1989
rect 49051 1961 49099 1989
rect 48789 -80 49099 1961
rect 48789 -108 48837 -80
rect 48865 -108 48899 -80
rect 48927 -108 48961 -80
rect 48989 -108 49023 -80
rect 49051 -108 49099 -80
rect 48789 -142 49099 -108
rect 48789 -170 48837 -142
rect 48865 -170 48899 -142
rect 48927 -170 48961 -142
rect 48989 -170 49023 -142
rect 49051 -170 49099 -142
rect 48789 -204 49099 -170
rect 48789 -232 48837 -204
rect 48865 -232 48899 -204
rect 48927 -232 48961 -204
rect 48989 -232 49023 -204
rect 49051 -232 49099 -204
rect 48789 -266 49099 -232
rect 48789 -294 48837 -266
rect 48865 -294 48899 -266
rect 48927 -294 48961 -266
rect 48989 -294 49023 -266
rect 49051 -294 49099 -266
rect 48789 -822 49099 -294
rect 50649 68175 50959 74345
rect 50649 68147 50697 68175
rect 50725 68147 50759 68175
rect 50787 68147 50821 68175
rect 50849 68147 50883 68175
rect 50911 68147 50959 68175
rect 50649 68113 50959 68147
rect 50649 68085 50697 68113
rect 50725 68085 50759 68113
rect 50787 68085 50821 68113
rect 50849 68085 50883 68113
rect 50911 68085 50959 68113
rect 50649 68051 50959 68085
rect 50649 68023 50697 68051
rect 50725 68023 50759 68051
rect 50787 68023 50821 68051
rect 50849 68023 50883 68051
rect 50911 68023 50959 68051
rect 50649 67989 50959 68023
rect 50649 67961 50697 67989
rect 50725 67961 50759 67989
rect 50787 67961 50821 67989
rect 50849 67961 50883 67989
rect 50911 67961 50959 67989
rect 50649 59175 50959 67961
rect 50649 59147 50697 59175
rect 50725 59147 50759 59175
rect 50787 59147 50821 59175
rect 50849 59147 50883 59175
rect 50911 59147 50959 59175
rect 50649 59113 50959 59147
rect 50649 59085 50697 59113
rect 50725 59085 50759 59113
rect 50787 59085 50821 59113
rect 50849 59085 50883 59113
rect 50911 59085 50959 59113
rect 50649 59051 50959 59085
rect 50649 59023 50697 59051
rect 50725 59023 50759 59051
rect 50787 59023 50821 59051
rect 50849 59023 50883 59051
rect 50911 59023 50959 59051
rect 50649 58989 50959 59023
rect 50649 58961 50697 58989
rect 50725 58961 50759 58989
rect 50787 58961 50821 58989
rect 50849 58961 50883 58989
rect 50911 58961 50959 58989
rect 50649 50175 50959 58961
rect 50649 50147 50697 50175
rect 50725 50147 50759 50175
rect 50787 50147 50821 50175
rect 50849 50147 50883 50175
rect 50911 50147 50959 50175
rect 50649 50113 50959 50147
rect 50649 50085 50697 50113
rect 50725 50085 50759 50113
rect 50787 50085 50821 50113
rect 50849 50085 50883 50113
rect 50911 50085 50959 50113
rect 50649 50051 50959 50085
rect 50649 50023 50697 50051
rect 50725 50023 50759 50051
rect 50787 50023 50821 50051
rect 50849 50023 50883 50051
rect 50911 50023 50959 50051
rect 50649 49989 50959 50023
rect 50649 49961 50697 49989
rect 50725 49961 50759 49989
rect 50787 49961 50821 49989
rect 50849 49961 50883 49989
rect 50911 49961 50959 49989
rect 50649 41175 50959 49961
rect 50649 41147 50697 41175
rect 50725 41147 50759 41175
rect 50787 41147 50821 41175
rect 50849 41147 50883 41175
rect 50911 41147 50959 41175
rect 50649 41113 50959 41147
rect 50649 41085 50697 41113
rect 50725 41085 50759 41113
rect 50787 41085 50821 41113
rect 50849 41085 50883 41113
rect 50911 41085 50959 41113
rect 50649 41051 50959 41085
rect 50649 41023 50697 41051
rect 50725 41023 50759 41051
rect 50787 41023 50821 41051
rect 50849 41023 50883 41051
rect 50911 41023 50959 41051
rect 50649 40989 50959 41023
rect 50649 40961 50697 40989
rect 50725 40961 50759 40989
rect 50787 40961 50821 40989
rect 50849 40961 50883 40989
rect 50911 40961 50959 40989
rect 50649 32175 50959 40961
rect 50649 32147 50697 32175
rect 50725 32147 50759 32175
rect 50787 32147 50821 32175
rect 50849 32147 50883 32175
rect 50911 32147 50959 32175
rect 50649 32113 50959 32147
rect 50649 32085 50697 32113
rect 50725 32085 50759 32113
rect 50787 32085 50821 32113
rect 50849 32085 50883 32113
rect 50911 32085 50959 32113
rect 50649 32051 50959 32085
rect 50649 32023 50697 32051
rect 50725 32023 50759 32051
rect 50787 32023 50821 32051
rect 50849 32023 50883 32051
rect 50911 32023 50959 32051
rect 50649 31989 50959 32023
rect 50649 31961 50697 31989
rect 50725 31961 50759 31989
rect 50787 31961 50821 31989
rect 50849 31961 50883 31989
rect 50911 31961 50959 31989
rect 50649 23175 50959 31961
rect 50649 23147 50697 23175
rect 50725 23147 50759 23175
rect 50787 23147 50821 23175
rect 50849 23147 50883 23175
rect 50911 23147 50959 23175
rect 50649 23113 50959 23147
rect 50649 23085 50697 23113
rect 50725 23085 50759 23113
rect 50787 23085 50821 23113
rect 50849 23085 50883 23113
rect 50911 23085 50959 23113
rect 50649 23051 50959 23085
rect 50649 23023 50697 23051
rect 50725 23023 50759 23051
rect 50787 23023 50821 23051
rect 50849 23023 50883 23051
rect 50911 23023 50959 23051
rect 50649 22989 50959 23023
rect 50649 22961 50697 22989
rect 50725 22961 50759 22989
rect 50787 22961 50821 22989
rect 50849 22961 50883 22989
rect 50911 22961 50959 22989
rect 50649 14175 50959 22961
rect 50649 14147 50697 14175
rect 50725 14147 50759 14175
rect 50787 14147 50821 14175
rect 50849 14147 50883 14175
rect 50911 14147 50959 14175
rect 50649 14113 50959 14147
rect 50649 14085 50697 14113
rect 50725 14085 50759 14113
rect 50787 14085 50821 14113
rect 50849 14085 50883 14113
rect 50911 14085 50959 14113
rect 50649 14051 50959 14085
rect 50649 14023 50697 14051
rect 50725 14023 50759 14051
rect 50787 14023 50821 14051
rect 50849 14023 50883 14051
rect 50911 14023 50959 14051
rect 50649 13989 50959 14023
rect 50649 13961 50697 13989
rect 50725 13961 50759 13989
rect 50787 13961 50821 13989
rect 50849 13961 50883 13989
rect 50911 13961 50959 13989
rect 50649 5175 50959 13961
rect 50649 5147 50697 5175
rect 50725 5147 50759 5175
rect 50787 5147 50821 5175
rect 50849 5147 50883 5175
rect 50911 5147 50959 5175
rect 50649 5113 50959 5147
rect 50649 5085 50697 5113
rect 50725 5085 50759 5113
rect 50787 5085 50821 5113
rect 50849 5085 50883 5113
rect 50911 5085 50959 5113
rect 50649 5051 50959 5085
rect 50649 5023 50697 5051
rect 50725 5023 50759 5051
rect 50787 5023 50821 5051
rect 50849 5023 50883 5051
rect 50911 5023 50959 5051
rect 50649 4989 50959 5023
rect 50649 4961 50697 4989
rect 50725 4961 50759 4989
rect 50787 4961 50821 4989
rect 50849 4961 50883 4989
rect 50911 4961 50959 4989
rect 50649 -560 50959 4961
rect 50649 -588 50697 -560
rect 50725 -588 50759 -560
rect 50787 -588 50821 -560
rect 50849 -588 50883 -560
rect 50911 -588 50959 -560
rect 50649 -622 50959 -588
rect 50649 -650 50697 -622
rect 50725 -650 50759 -622
rect 50787 -650 50821 -622
rect 50849 -650 50883 -622
rect 50911 -650 50959 -622
rect 50649 -684 50959 -650
rect 50649 -712 50697 -684
rect 50725 -712 50759 -684
rect 50787 -712 50821 -684
rect 50849 -712 50883 -684
rect 50911 -712 50959 -684
rect 50649 -746 50959 -712
rect 50649 -774 50697 -746
rect 50725 -774 50759 -746
rect 50787 -774 50821 -746
rect 50849 -774 50883 -746
rect 50911 -774 50959 -746
rect 50649 -822 50959 -774
rect 64149 74175 64459 74345
rect 64149 74147 64197 74175
rect 64225 74147 64259 74175
rect 64287 74147 64321 74175
rect 64349 74147 64383 74175
rect 64411 74147 64459 74175
rect 64149 74113 64459 74147
rect 64149 74085 64197 74113
rect 64225 74085 64259 74113
rect 64287 74085 64321 74113
rect 64349 74085 64383 74113
rect 64411 74085 64459 74113
rect 64149 74051 64459 74085
rect 64149 74023 64197 74051
rect 64225 74023 64259 74051
rect 64287 74023 64321 74051
rect 64349 74023 64383 74051
rect 64411 74023 64459 74051
rect 64149 73989 64459 74023
rect 64149 73961 64197 73989
rect 64225 73961 64259 73989
rect 64287 73961 64321 73989
rect 64349 73961 64383 73989
rect 64411 73961 64459 73989
rect 64149 65175 64459 73961
rect 64149 65147 64197 65175
rect 64225 65147 64259 65175
rect 64287 65147 64321 65175
rect 64349 65147 64383 65175
rect 64411 65147 64459 65175
rect 64149 65113 64459 65147
rect 64149 65085 64197 65113
rect 64225 65085 64259 65113
rect 64287 65085 64321 65113
rect 64349 65085 64383 65113
rect 64411 65085 64459 65113
rect 64149 65051 64459 65085
rect 64149 65023 64197 65051
rect 64225 65023 64259 65051
rect 64287 65023 64321 65051
rect 64349 65023 64383 65051
rect 64411 65023 64459 65051
rect 64149 64989 64459 65023
rect 64149 64961 64197 64989
rect 64225 64961 64259 64989
rect 64287 64961 64321 64989
rect 64349 64961 64383 64989
rect 64411 64961 64459 64989
rect 64149 56175 64459 64961
rect 64149 56147 64197 56175
rect 64225 56147 64259 56175
rect 64287 56147 64321 56175
rect 64349 56147 64383 56175
rect 64411 56147 64459 56175
rect 64149 56113 64459 56147
rect 64149 56085 64197 56113
rect 64225 56085 64259 56113
rect 64287 56085 64321 56113
rect 64349 56085 64383 56113
rect 64411 56085 64459 56113
rect 64149 56051 64459 56085
rect 64149 56023 64197 56051
rect 64225 56023 64259 56051
rect 64287 56023 64321 56051
rect 64349 56023 64383 56051
rect 64411 56023 64459 56051
rect 64149 55989 64459 56023
rect 64149 55961 64197 55989
rect 64225 55961 64259 55989
rect 64287 55961 64321 55989
rect 64349 55961 64383 55989
rect 64411 55961 64459 55989
rect 64149 47175 64459 55961
rect 64149 47147 64197 47175
rect 64225 47147 64259 47175
rect 64287 47147 64321 47175
rect 64349 47147 64383 47175
rect 64411 47147 64459 47175
rect 64149 47113 64459 47147
rect 64149 47085 64197 47113
rect 64225 47085 64259 47113
rect 64287 47085 64321 47113
rect 64349 47085 64383 47113
rect 64411 47085 64459 47113
rect 64149 47051 64459 47085
rect 64149 47023 64197 47051
rect 64225 47023 64259 47051
rect 64287 47023 64321 47051
rect 64349 47023 64383 47051
rect 64411 47023 64459 47051
rect 64149 46989 64459 47023
rect 64149 46961 64197 46989
rect 64225 46961 64259 46989
rect 64287 46961 64321 46989
rect 64349 46961 64383 46989
rect 64411 46961 64459 46989
rect 64149 38175 64459 46961
rect 64149 38147 64197 38175
rect 64225 38147 64259 38175
rect 64287 38147 64321 38175
rect 64349 38147 64383 38175
rect 64411 38147 64459 38175
rect 64149 38113 64459 38147
rect 64149 38085 64197 38113
rect 64225 38085 64259 38113
rect 64287 38085 64321 38113
rect 64349 38085 64383 38113
rect 64411 38085 64459 38113
rect 64149 38051 64459 38085
rect 64149 38023 64197 38051
rect 64225 38023 64259 38051
rect 64287 38023 64321 38051
rect 64349 38023 64383 38051
rect 64411 38023 64459 38051
rect 64149 37989 64459 38023
rect 64149 37961 64197 37989
rect 64225 37961 64259 37989
rect 64287 37961 64321 37989
rect 64349 37961 64383 37989
rect 64411 37961 64459 37989
rect 64149 29175 64459 37961
rect 64149 29147 64197 29175
rect 64225 29147 64259 29175
rect 64287 29147 64321 29175
rect 64349 29147 64383 29175
rect 64411 29147 64459 29175
rect 64149 29113 64459 29147
rect 64149 29085 64197 29113
rect 64225 29085 64259 29113
rect 64287 29085 64321 29113
rect 64349 29085 64383 29113
rect 64411 29085 64459 29113
rect 64149 29051 64459 29085
rect 64149 29023 64197 29051
rect 64225 29023 64259 29051
rect 64287 29023 64321 29051
rect 64349 29023 64383 29051
rect 64411 29023 64459 29051
rect 64149 28989 64459 29023
rect 64149 28961 64197 28989
rect 64225 28961 64259 28989
rect 64287 28961 64321 28989
rect 64349 28961 64383 28989
rect 64411 28961 64459 28989
rect 64149 20175 64459 28961
rect 64149 20147 64197 20175
rect 64225 20147 64259 20175
rect 64287 20147 64321 20175
rect 64349 20147 64383 20175
rect 64411 20147 64459 20175
rect 64149 20113 64459 20147
rect 64149 20085 64197 20113
rect 64225 20085 64259 20113
rect 64287 20085 64321 20113
rect 64349 20085 64383 20113
rect 64411 20085 64459 20113
rect 64149 20051 64459 20085
rect 64149 20023 64197 20051
rect 64225 20023 64259 20051
rect 64287 20023 64321 20051
rect 64349 20023 64383 20051
rect 64411 20023 64459 20051
rect 64149 19989 64459 20023
rect 64149 19961 64197 19989
rect 64225 19961 64259 19989
rect 64287 19961 64321 19989
rect 64349 19961 64383 19989
rect 64411 19961 64459 19989
rect 64149 11175 64459 19961
rect 64149 11147 64197 11175
rect 64225 11147 64259 11175
rect 64287 11147 64321 11175
rect 64349 11147 64383 11175
rect 64411 11147 64459 11175
rect 64149 11113 64459 11147
rect 64149 11085 64197 11113
rect 64225 11085 64259 11113
rect 64287 11085 64321 11113
rect 64349 11085 64383 11113
rect 64411 11085 64459 11113
rect 64149 11051 64459 11085
rect 64149 11023 64197 11051
rect 64225 11023 64259 11051
rect 64287 11023 64321 11051
rect 64349 11023 64383 11051
rect 64411 11023 64459 11051
rect 64149 10989 64459 11023
rect 64149 10961 64197 10989
rect 64225 10961 64259 10989
rect 64287 10961 64321 10989
rect 64349 10961 64383 10989
rect 64411 10961 64459 10989
rect 64149 2175 64459 10961
rect 64149 2147 64197 2175
rect 64225 2147 64259 2175
rect 64287 2147 64321 2175
rect 64349 2147 64383 2175
rect 64411 2147 64459 2175
rect 64149 2113 64459 2147
rect 64149 2085 64197 2113
rect 64225 2085 64259 2113
rect 64287 2085 64321 2113
rect 64349 2085 64383 2113
rect 64411 2085 64459 2113
rect 64149 2051 64459 2085
rect 64149 2023 64197 2051
rect 64225 2023 64259 2051
rect 64287 2023 64321 2051
rect 64349 2023 64383 2051
rect 64411 2023 64459 2051
rect 64149 1989 64459 2023
rect 64149 1961 64197 1989
rect 64225 1961 64259 1989
rect 64287 1961 64321 1989
rect 64349 1961 64383 1989
rect 64411 1961 64459 1989
rect 64149 -80 64459 1961
rect 64149 -108 64197 -80
rect 64225 -108 64259 -80
rect 64287 -108 64321 -80
rect 64349 -108 64383 -80
rect 64411 -108 64459 -80
rect 64149 -142 64459 -108
rect 64149 -170 64197 -142
rect 64225 -170 64259 -142
rect 64287 -170 64321 -142
rect 64349 -170 64383 -142
rect 64411 -170 64459 -142
rect 64149 -204 64459 -170
rect 64149 -232 64197 -204
rect 64225 -232 64259 -204
rect 64287 -232 64321 -204
rect 64349 -232 64383 -204
rect 64411 -232 64459 -204
rect 64149 -266 64459 -232
rect 64149 -294 64197 -266
rect 64225 -294 64259 -266
rect 64287 -294 64321 -266
rect 64349 -294 64383 -266
rect 64411 -294 64459 -266
rect 64149 -822 64459 -294
rect 66009 68175 66319 74345
rect 66009 68147 66057 68175
rect 66085 68147 66119 68175
rect 66147 68147 66181 68175
rect 66209 68147 66243 68175
rect 66271 68147 66319 68175
rect 66009 68113 66319 68147
rect 66009 68085 66057 68113
rect 66085 68085 66119 68113
rect 66147 68085 66181 68113
rect 66209 68085 66243 68113
rect 66271 68085 66319 68113
rect 66009 68051 66319 68085
rect 66009 68023 66057 68051
rect 66085 68023 66119 68051
rect 66147 68023 66181 68051
rect 66209 68023 66243 68051
rect 66271 68023 66319 68051
rect 66009 67989 66319 68023
rect 66009 67961 66057 67989
rect 66085 67961 66119 67989
rect 66147 67961 66181 67989
rect 66209 67961 66243 67989
rect 66271 67961 66319 67989
rect 66009 59175 66319 67961
rect 66009 59147 66057 59175
rect 66085 59147 66119 59175
rect 66147 59147 66181 59175
rect 66209 59147 66243 59175
rect 66271 59147 66319 59175
rect 66009 59113 66319 59147
rect 66009 59085 66057 59113
rect 66085 59085 66119 59113
rect 66147 59085 66181 59113
rect 66209 59085 66243 59113
rect 66271 59085 66319 59113
rect 66009 59051 66319 59085
rect 66009 59023 66057 59051
rect 66085 59023 66119 59051
rect 66147 59023 66181 59051
rect 66209 59023 66243 59051
rect 66271 59023 66319 59051
rect 66009 58989 66319 59023
rect 66009 58961 66057 58989
rect 66085 58961 66119 58989
rect 66147 58961 66181 58989
rect 66209 58961 66243 58989
rect 66271 58961 66319 58989
rect 66009 50175 66319 58961
rect 66009 50147 66057 50175
rect 66085 50147 66119 50175
rect 66147 50147 66181 50175
rect 66209 50147 66243 50175
rect 66271 50147 66319 50175
rect 66009 50113 66319 50147
rect 66009 50085 66057 50113
rect 66085 50085 66119 50113
rect 66147 50085 66181 50113
rect 66209 50085 66243 50113
rect 66271 50085 66319 50113
rect 66009 50051 66319 50085
rect 66009 50023 66057 50051
rect 66085 50023 66119 50051
rect 66147 50023 66181 50051
rect 66209 50023 66243 50051
rect 66271 50023 66319 50051
rect 66009 49989 66319 50023
rect 66009 49961 66057 49989
rect 66085 49961 66119 49989
rect 66147 49961 66181 49989
rect 66209 49961 66243 49989
rect 66271 49961 66319 49989
rect 66009 41175 66319 49961
rect 66009 41147 66057 41175
rect 66085 41147 66119 41175
rect 66147 41147 66181 41175
rect 66209 41147 66243 41175
rect 66271 41147 66319 41175
rect 66009 41113 66319 41147
rect 66009 41085 66057 41113
rect 66085 41085 66119 41113
rect 66147 41085 66181 41113
rect 66209 41085 66243 41113
rect 66271 41085 66319 41113
rect 66009 41051 66319 41085
rect 66009 41023 66057 41051
rect 66085 41023 66119 41051
rect 66147 41023 66181 41051
rect 66209 41023 66243 41051
rect 66271 41023 66319 41051
rect 66009 40989 66319 41023
rect 66009 40961 66057 40989
rect 66085 40961 66119 40989
rect 66147 40961 66181 40989
rect 66209 40961 66243 40989
rect 66271 40961 66319 40989
rect 66009 32175 66319 40961
rect 66009 32147 66057 32175
rect 66085 32147 66119 32175
rect 66147 32147 66181 32175
rect 66209 32147 66243 32175
rect 66271 32147 66319 32175
rect 66009 32113 66319 32147
rect 66009 32085 66057 32113
rect 66085 32085 66119 32113
rect 66147 32085 66181 32113
rect 66209 32085 66243 32113
rect 66271 32085 66319 32113
rect 66009 32051 66319 32085
rect 66009 32023 66057 32051
rect 66085 32023 66119 32051
rect 66147 32023 66181 32051
rect 66209 32023 66243 32051
rect 66271 32023 66319 32051
rect 66009 31989 66319 32023
rect 66009 31961 66057 31989
rect 66085 31961 66119 31989
rect 66147 31961 66181 31989
rect 66209 31961 66243 31989
rect 66271 31961 66319 31989
rect 66009 23175 66319 31961
rect 66009 23147 66057 23175
rect 66085 23147 66119 23175
rect 66147 23147 66181 23175
rect 66209 23147 66243 23175
rect 66271 23147 66319 23175
rect 66009 23113 66319 23147
rect 66009 23085 66057 23113
rect 66085 23085 66119 23113
rect 66147 23085 66181 23113
rect 66209 23085 66243 23113
rect 66271 23085 66319 23113
rect 66009 23051 66319 23085
rect 66009 23023 66057 23051
rect 66085 23023 66119 23051
rect 66147 23023 66181 23051
rect 66209 23023 66243 23051
rect 66271 23023 66319 23051
rect 66009 22989 66319 23023
rect 66009 22961 66057 22989
rect 66085 22961 66119 22989
rect 66147 22961 66181 22989
rect 66209 22961 66243 22989
rect 66271 22961 66319 22989
rect 66009 14175 66319 22961
rect 66009 14147 66057 14175
rect 66085 14147 66119 14175
rect 66147 14147 66181 14175
rect 66209 14147 66243 14175
rect 66271 14147 66319 14175
rect 66009 14113 66319 14147
rect 66009 14085 66057 14113
rect 66085 14085 66119 14113
rect 66147 14085 66181 14113
rect 66209 14085 66243 14113
rect 66271 14085 66319 14113
rect 66009 14051 66319 14085
rect 66009 14023 66057 14051
rect 66085 14023 66119 14051
rect 66147 14023 66181 14051
rect 66209 14023 66243 14051
rect 66271 14023 66319 14051
rect 66009 13989 66319 14023
rect 66009 13961 66057 13989
rect 66085 13961 66119 13989
rect 66147 13961 66181 13989
rect 66209 13961 66243 13989
rect 66271 13961 66319 13989
rect 66009 5175 66319 13961
rect 66009 5147 66057 5175
rect 66085 5147 66119 5175
rect 66147 5147 66181 5175
rect 66209 5147 66243 5175
rect 66271 5147 66319 5175
rect 66009 5113 66319 5147
rect 66009 5085 66057 5113
rect 66085 5085 66119 5113
rect 66147 5085 66181 5113
rect 66209 5085 66243 5113
rect 66271 5085 66319 5113
rect 66009 5051 66319 5085
rect 66009 5023 66057 5051
rect 66085 5023 66119 5051
rect 66147 5023 66181 5051
rect 66209 5023 66243 5051
rect 66271 5023 66319 5051
rect 66009 4989 66319 5023
rect 66009 4961 66057 4989
rect 66085 4961 66119 4989
rect 66147 4961 66181 4989
rect 66209 4961 66243 4989
rect 66271 4961 66319 4989
rect 66009 -560 66319 4961
rect 66009 -588 66057 -560
rect 66085 -588 66119 -560
rect 66147 -588 66181 -560
rect 66209 -588 66243 -560
rect 66271 -588 66319 -560
rect 66009 -622 66319 -588
rect 66009 -650 66057 -622
rect 66085 -650 66119 -622
rect 66147 -650 66181 -622
rect 66209 -650 66243 -622
rect 66271 -650 66319 -622
rect 66009 -684 66319 -650
rect 66009 -712 66057 -684
rect 66085 -712 66119 -684
rect 66147 -712 66181 -684
rect 66209 -712 66243 -684
rect 66271 -712 66319 -684
rect 66009 -746 66319 -712
rect 66009 -774 66057 -746
rect 66085 -774 66119 -746
rect 66147 -774 66181 -746
rect 66209 -774 66243 -746
rect 66271 -774 66319 -746
rect 66009 -822 66319 -774
rect 79509 74175 79819 82961
rect 79509 74147 79557 74175
rect 79585 74147 79619 74175
rect 79647 74147 79681 74175
rect 79709 74147 79743 74175
rect 79771 74147 79819 74175
rect 79509 74113 79819 74147
rect 79509 74085 79557 74113
rect 79585 74085 79619 74113
rect 79647 74085 79681 74113
rect 79709 74085 79743 74113
rect 79771 74085 79819 74113
rect 79509 74051 79819 74085
rect 79509 74023 79557 74051
rect 79585 74023 79619 74051
rect 79647 74023 79681 74051
rect 79709 74023 79743 74051
rect 79771 74023 79819 74051
rect 79509 73989 79819 74023
rect 79509 73961 79557 73989
rect 79585 73961 79619 73989
rect 79647 73961 79681 73989
rect 79709 73961 79743 73989
rect 79771 73961 79819 73989
rect 79509 65175 79819 73961
rect 79509 65147 79557 65175
rect 79585 65147 79619 65175
rect 79647 65147 79681 65175
rect 79709 65147 79743 65175
rect 79771 65147 79819 65175
rect 79509 65113 79819 65147
rect 79509 65085 79557 65113
rect 79585 65085 79619 65113
rect 79647 65085 79681 65113
rect 79709 65085 79743 65113
rect 79771 65085 79819 65113
rect 79509 65051 79819 65085
rect 79509 65023 79557 65051
rect 79585 65023 79619 65051
rect 79647 65023 79681 65051
rect 79709 65023 79743 65051
rect 79771 65023 79819 65051
rect 79509 64989 79819 65023
rect 79509 64961 79557 64989
rect 79585 64961 79619 64989
rect 79647 64961 79681 64989
rect 79709 64961 79743 64989
rect 79771 64961 79819 64989
rect 79509 56175 79819 64961
rect 79509 56147 79557 56175
rect 79585 56147 79619 56175
rect 79647 56147 79681 56175
rect 79709 56147 79743 56175
rect 79771 56147 79819 56175
rect 79509 56113 79819 56147
rect 79509 56085 79557 56113
rect 79585 56085 79619 56113
rect 79647 56085 79681 56113
rect 79709 56085 79743 56113
rect 79771 56085 79819 56113
rect 79509 56051 79819 56085
rect 79509 56023 79557 56051
rect 79585 56023 79619 56051
rect 79647 56023 79681 56051
rect 79709 56023 79743 56051
rect 79771 56023 79819 56051
rect 79509 55989 79819 56023
rect 79509 55961 79557 55989
rect 79585 55961 79619 55989
rect 79647 55961 79681 55989
rect 79709 55961 79743 55989
rect 79771 55961 79819 55989
rect 79509 47175 79819 55961
rect 79509 47147 79557 47175
rect 79585 47147 79619 47175
rect 79647 47147 79681 47175
rect 79709 47147 79743 47175
rect 79771 47147 79819 47175
rect 79509 47113 79819 47147
rect 79509 47085 79557 47113
rect 79585 47085 79619 47113
rect 79647 47085 79681 47113
rect 79709 47085 79743 47113
rect 79771 47085 79819 47113
rect 79509 47051 79819 47085
rect 79509 47023 79557 47051
rect 79585 47023 79619 47051
rect 79647 47023 79681 47051
rect 79709 47023 79743 47051
rect 79771 47023 79819 47051
rect 79509 46989 79819 47023
rect 79509 46961 79557 46989
rect 79585 46961 79619 46989
rect 79647 46961 79681 46989
rect 79709 46961 79743 46989
rect 79771 46961 79819 46989
rect 79509 38175 79819 46961
rect 79509 38147 79557 38175
rect 79585 38147 79619 38175
rect 79647 38147 79681 38175
rect 79709 38147 79743 38175
rect 79771 38147 79819 38175
rect 79509 38113 79819 38147
rect 79509 38085 79557 38113
rect 79585 38085 79619 38113
rect 79647 38085 79681 38113
rect 79709 38085 79743 38113
rect 79771 38085 79819 38113
rect 79509 38051 79819 38085
rect 79509 38023 79557 38051
rect 79585 38023 79619 38051
rect 79647 38023 79681 38051
rect 79709 38023 79743 38051
rect 79771 38023 79819 38051
rect 79509 37989 79819 38023
rect 79509 37961 79557 37989
rect 79585 37961 79619 37989
rect 79647 37961 79681 37989
rect 79709 37961 79743 37989
rect 79771 37961 79819 37989
rect 79509 29175 79819 37961
rect 79509 29147 79557 29175
rect 79585 29147 79619 29175
rect 79647 29147 79681 29175
rect 79709 29147 79743 29175
rect 79771 29147 79819 29175
rect 79509 29113 79819 29147
rect 79509 29085 79557 29113
rect 79585 29085 79619 29113
rect 79647 29085 79681 29113
rect 79709 29085 79743 29113
rect 79771 29085 79819 29113
rect 79509 29051 79819 29085
rect 79509 29023 79557 29051
rect 79585 29023 79619 29051
rect 79647 29023 79681 29051
rect 79709 29023 79743 29051
rect 79771 29023 79819 29051
rect 79509 28989 79819 29023
rect 79509 28961 79557 28989
rect 79585 28961 79619 28989
rect 79647 28961 79681 28989
rect 79709 28961 79743 28989
rect 79771 28961 79819 28989
rect 79509 20175 79819 28961
rect 79509 20147 79557 20175
rect 79585 20147 79619 20175
rect 79647 20147 79681 20175
rect 79709 20147 79743 20175
rect 79771 20147 79819 20175
rect 79509 20113 79819 20147
rect 79509 20085 79557 20113
rect 79585 20085 79619 20113
rect 79647 20085 79681 20113
rect 79709 20085 79743 20113
rect 79771 20085 79819 20113
rect 79509 20051 79819 20085
rect 79509 20023 79557 20051
rect 79585 20023 79619 20051
rect 79647 20023 79681 20051
rect 79709 20023 79743 20051
rect 79771 20023 79819 20051
rect 79509 19989 79819 20023
rect 79509 19961 79557 19989
rect 79585 19961 79619 19989
rect 79647 19961 79681 19989
rect 79709 19961 79743 19989
rect 79771 19961 79819 19989
rect 79509 11175 79819 19961
rect 79509 11147 79557 11175
rect 79585 11147 79619 11175
rect 79647 11147 79681 11175
rect 79709 11147 79743 11175
rect 79771 11147 79819 11175
rect 79509 11113 79819 11147
rect 79509 11085 79557 11113
rect 79585 11085 79619 11113
rect 79647 11085 79681 11113
rect 79709 11085 79743 11113
rect 79771 11085 79819 11113
rect 79509 11051 79819 11085
rect 79509 11023 79557 11051
rect 79585 11023 79619 11051
rect 79647 11023 79681 11051
rect 79709 11023 79743 11051
rect 79771 11023 79819 11051
rect 79509 10989 79819 11023
rect 79509 10961 79557 10989
rect 79585 10961 79619 10989
rect 79647 10961 79681 10989
rect 79709 10961 79743 10989
rect 79771 10961 79819 10989
rect 79509 2175 79819 10961
rect 79509 2147 79557 2175
rect 79585 2147 79619 2175
rect 79647 2147 79681 2175
rect 79709 2147 79743 2175
rect 79771 2147 79819 2175
rect 79509 2113 79819 2147
rect 79509 2085 79557 2113
rect 79585 2085 79619 2113
rect 79647 2085 79681 2113
rect 79709 2085 79743 2113
rect 79771 2085 79819 2113
rect 79509 2051 79819 2085
rect 79509 2023 79557 2051
rect 79585 2023 79619 2051
rect 79647 2023 79681 2051
rect 79709 2023 79743 2051
rect 79771 2023 79819 2051
rect 79509 1989 79819 2023
rect 79509 1961 79557 1989
rect 79585 1961 79619 1989
rect 79647 1961 79681 1989
rect 79709 1961 79743 1989
rect 79771 1961 79819 1989
rect 79509 -80 79819 1961
rect 79509 -108 79557 -80
rect 79585 -108 79619 -80
rect 79647 -108 79681 -80
rect 79709 -108 79743 -80
rect 79771 -108 79819 -80
rect 79509 -142 79819 -108
rect 79509 -170 79557 -142
rect 79585 -170 79619 -142
rect 79647 -170 79681 -142
rect 79709 -170 79743 -142
rect 79771 -170 79819 -142
rect 79509 -204 79819 -170
rect 79509 -232 79557 -204
rect 79585 -232 79619 -204
rect 79647 -232 79681 -204
rect 79709 -232 79743 -204
rect 79771 -232 79819 -204
rect 79509 -266 79819 -232
rect 79509 -294 79557 -266
rect 79585 -294 79619 -266
rect 79647 -294 79681 -266
rect 79709 -294 79743 -266
rect 79771 -294 79819 -266
rect 79509 -822 79819 -294
rect 81369 167175 81679 170745
rect 81369 167147 81417 167175
rect 81445 167147 81479 167175
rect 81507 167147 81541 167175
rect 81569 167147 81603 167175
rect 81631 167147 81679 167175
rect 81369 167113 81679 167147
rect 81369 167085 81417 167113
rect 81445 167085 81479 167113
rect 81507 167085 81541 167113
rect 81569 167085 81603 167113
rect 81631 167085 81679 167113
rect 81369 167051 81679 167085
rect 81369 167023 81417 167051
rect 81445 167023 81479 167051
rect 81507 167023 81541 167051
rect 81569 167023 81603 167051
rect 81631 167023 81679 167051
rect 81369 166989 81679 167023
rect 81369 166961 81417 166989
rect 81445 166961 81479 166989
rect 81507 166961 81541 166989
rect 81569 166961 81603 166989
rect 81631 166961 81679 166989
rect 81369 158175 81679 166961
rect 94869 164175 95179 172961
rect 94869 164147 94917 164175
rect 94945 164147 94979 164175
rect 95007 164147 95041 164175
rect 95069 164147 95103 164175
rect 95131 164147 95179 164175
rect 94869 164113 95179 164147
rect 94869 164085 94917 164113
rect 94945 164085 94979 164113
rect 95007 164085 95041 164113
rect 95069 164085 95103 164113
rect 95131 164085 95179 164113
rect 94869 164051 95179 164085
rect 94869 164023 94917 164051
rect 94945 164023 94979 164051
rect 95007 164023 95041 164051
rect 95069 164023 95103 164051
rect 95131 164023 95179 164051
rect 94869 163989 95179 164023
rect 94869 163961 94917 163989
rect 94945 163961 94979 163989
rect 95007 163961 95041 163989
rect 95069 163961 95103 163989
rect 95131 163961 95179 163989
rect 81369 158147 81417 158175
rect 81445 158147 81479 158175
rect 81507 158147 81541 158175
rect 81569 158147 81603 158175
rect 81631 158147 81679 158175
rect 81369 158113 81679 158147
rect 81369 158085 81417 158113
rect 81445 158085 81479 158113
rect 81507 158085 81541 158113
rect 81569 158085 81603 158113
rect 81631 158085 81679 158113
rect 81369 158051 81679 158085
rect 81369 158023 81417 158051
rect 81445 158023 81479 158051
rect 81507 158023 81541 158051
rect 81569 158023 81603 158051
rect 81631 158023 81679 158051
rect 81369 157989 81679 158023
rect 81369 157961 81417 157989
rect 81445 157961 81479 157989
rect 81507 157961 81541 157989
rect 81569 157961 81603 157989
rect 81631 157961 81679 157989
rect 81369 149175 81679 157961
rect 85984 158175 86144 158192
rect 85984 158147 86019 158175
rect 86047 158147 86081 158175
rect 86109 158147 86144 158175
rect 85984 158113 86144 158147
rect 85984 158085 86019 158113
rect 86047 158085 86081 158113
rect 86109 158085 86144 158113
rect 85984 158051 86144 158085
rect 85984 158023 86019 158051
rect 86047 158023 86081 158051
rect 86109 158023 86144 158051
rect 85984 157989 86144 158023
rect 85984 157961 86019 157989
rect 86047 157961 86081 157989
rect 86109 157961 86144 157989
rect 85984 157944 86144 157961
rect 93664 155175 93824 155192
rect 93664 155147 93699 155175
rect 93727 155147 93761 155175
rect 93789 155147 93824 155175
rect 93664 155113 93824 155147
rect 93664 155085 93699 155113
rect 93727 155085 93761 155113
rect 93789 155085 93824 155113
rect 93664 155051 93824 155085
rect 93664 155023 93699 155051
rect 93727 155023 93761 155051
rect 93789 155023 93824 155051
rect 93664 154989 93824 155023
rect 93664 154961 93699 154989
rect 93727 154961 93761 154989
rect 93789 154961 93824 154989
rect 93664 154944 93824 154961
rect 94869 155175 95179 163961
rect 94869 155147 94917 155175
rect 94945 155147 94979 155175
rect 95007 155147 95041 155175
rect 95069 155147 95103 155175
rect 95131 155147 95179 155175
rect 94869 155113 95179 155147
rect 94869 155085 94917 155113
rect 94945 155085 94979 155113
rect 95007 155085 95041 155113
rect 95069 155085 95103 155113
rect 95131 155085 95179 155113
rect 94869 155051 95179 155085
rect 94869 155023 94917 155051
rect 94945 155023 94979 155051
rect 95007 155023 95041 155051
rect 95069 155023 95103 155051
rect 95131 155023 95179 155051
rect 94869 154989 95179 155023
rect 94869 154961 94917 154989
rect 94945 154961 94979 154989
rect 95007 154961 95041 154989
rect 95069 154961 95103 154989
rect 95131 154961 95179 154989
rect 81369 149147 81417 149175
rect 81445 149147 81479 149175
rect 81507 149147 81541 149175
rect 81569 149147 81603 149175
rect 81631 149147 81679 149175
rect 81369 149113 81679 149147
rect 81369 149085 81417 149113
rect 81445 149085 81479 149113
rect 81507 149085 81541 149113
rect 81569 149085 81603 149113
rect 81631 149085 81679 149113
rect 81369 149051 81679 149085
rect 81369 149023 81417 149051
rect 81445 149023 81479 149051
rect 81507 149023 81541 149051
rect 81569 149023 81603 149051
rect 81631 149023 81679 149051
rect 81369 148989 81679 149023
rect 81369 148961 81417 148989
rect 81445 148961 81479 148989
rect 81507 148961 81541 148989
rect 81569 148961 81603 148989
rect 81631 148961 81679 148989
rect 81369 140175 81679 148961
rect 85984 149175 86144 149192
rect 85984 149147 86019 149175
rect 86047 149147 86081 149175
rect 86109 149147 86144 149175
rect 85984 149113 86144 149147
rect 85984 149085 86019 149113
rect 86047 149085 86081 149113
rect 86109 149085 86144 149113
rect 85984 149051 86144 149085
rect 85984 149023 86019 149051
rect 86047 149023 86081 149051
rect 86109 149023 86144 149051
rect 85984 148989 86144 149023
rect 85984 148961 86019 148989
rect 86047 148961 86081 148989
rect 86109 148961 86144 148989
rect 85984 148944 86144 148961
rect 93664 146175 93824 146192
rect 93664 146147 93699 146175
rect 93727 146147 93761 146175
rect 93789 146147 93824 146175
rect 93664 146113 93824 146147
rect 93664 146085 93699 146113
rect 93727 146085 93761 146113
rect 93789 146085 93824 146113
rect 93664 146051 93824 146085
rect 93664 146023 93699 146051
rect 93727 146023 93761 146051
rect 93789 146023 93824 146051
rect 93664 145989 93824 146023
rect 93664 145961 93699 145989
rect 93727 145961 93761 145989
rect 93789 145961 93824 145989
rect 93664 145944 93824 145961
rect 94869 146175 95179 154961
rect 94869 146147 94917 146175
rect 94945 146147 94979 146175
rect 95007 146147 95041 146175
rect 95069 146147 95103 146175
rect 95131 146147 95179 146175
rect 94869 146113 95179 146147
rect 94869 146085 94917 146113
rect 94945 146085 94979 146113
rect 95007 146085 95041 146113
rect 95069 146085 95103 146113
rect 95131 146085 95179 146113
rect 94869 146051 95179 146085
rect 94869 146023 94917 146051
rect 94945 146023 94979 146051
rect 95007 146023 95041 146051
rect 95069 146023 95103 146051
rect 95131 146023 95179 146051
rect 94869 145989 95179 146023
rect 94869 145961 94917 145989
rect 94945 145961 94979 145989
rect 95007 145961 95041 145989
rect 95069 145961 95103 145989
rect 95131 145961 95179 145989
rect 81369 140147 81417 140175
rect 81445 140147 81479 140175
rect 81507 140147 81541 140175
rect 81569 140147 81603 140175
rect 81631 140147 81679 140175
rect 81369 140113 81679 140147
rect 81369 140085 81417 140113
rect 81445 140085 81479 140113
rect 81507 140085 81541 140113
rect 81569 140085 81603 140113
rect 81631 140085 81679 140113
rect 81369 140051 81679 140085
rect 81369 140023 81417 140051
rect 81445 140023 81479 140051
rect 81507 140023 81541 140051
rect 81569 140023 81603 140051
rect 81631 140023 81679 140051
rect 81369 139989 81679 140023
rect 81369 139961 81417 139989
rect 81445 139961 81479 139989
rect 81507 139961 81541 139989
rect 81569 139961 81603 139989
rect 81631 139961 81679 139989
rect 81369 131175 81679 139961
rect 85984 140175 86144 140192
rect 85984 140147 86019 140175
rect 86047 140147 86081 140175
rect 86109 140147 86144 140175
rect 85984 140113 86144 140147
rect 85984 140085 86019 140113
rect 86047 140085 86081 140113
rect 86109 140085 86144 140113
rect 85984 140051 86144 140085
rect 85984 140023 86019 140051
rect 86047 140023 86081 140051
rect 86109 140023 86144 140051
rect 85984 139989 86144 140023
rect 85984 139961 86019 139989
rect 86047 139961 86081 139989
rect 86109 139961 86144 139989
rect 85984 139944 86144 139961
rect 93664 137175 93824 137192
rect 93664 137147 93699 137175
rect 93727 137147 93761 137175
rect 93789 137147 93824 137175
rect 93664 137113 93824 137147
rect 93664 137085 93699 137113
rect 93727 137085 93761 137113
rect 93789 137085 93824 137113
rect 93664 137051 93824 137085
rect 93664 137023 93699 137051
rect 93727 137023 93761 137051
rect 93789 137023 93824 137051
rect 93664 136989 93824 137023
rect 93664 136961 93699 136989
rect 93727 136961 93761 136989
rect 93789 136961 93824 136989
rect 93664 136944 93824 136961
rect 94869 137175 95179 145961
rect 94869 137147 94917 137175
rect 94945 137147 94979 137175
rect 95007 137147 95041 137175
rect 95069 137147 95103 137175
rect 95131 137147 95179 137175
rect 94869 137113 95179 137147
rect 94869 137085 94917 137113
rect 94945 137085 94979 137113
rect 95007 137085 95041 137113
rect 95069 137085 95103 137113
rect 95131 137085 95179 137113
rect 94869 137051 95179 137085
rect 94869 137023 94917 137051
rect 94945 137023 94979 137051
rect 95007 137023 95041 137051
rect 95069 137023 95103 137051
rect 95131 137023 95179 137051
rect 94869 136989 95179 137023
rect 94869 136961 94917 136989
rect 94945 136961 94979 136989
rect 95007 136961 95041 136989
rect 95069 136961 95103 136989
rect 95131 136961 95179 136989
rect 81369 131147 81417 131175
rect 81445 131147 81479 131175
rect 81507 131147 81541 131175
rect 81569 131147 81603 131175
rect 81631 131147 81679 131175
rect 81369 131113 81679 131147
rect 81369 131085 81417 131113
rect 81445 131085 81479 131113
rect 81507 131085 81541 131113
rect 81569 131085 81603 131113
rect 81631 131085 81679 131113
rect 81369 131051 81679 131085
rect 81369 131023 81417 131051
rect 81445 131023 81479 131051
rect 81507 131023 81541 131051
rect 81569 131023 81603 131051
rect 81631 131023 81679 131051
rect 81369 130989 81679 131023
rect 81369 130961 81417 130989
rect 81445 130961 81479 130989
rect 81507 130961 81541 130989
rect 81569 130961 81603 130989
rect 81631 130961 81679 130989
rect 81369 122175 81679 130961
rect 81369 122147 81417 122175
rect 81445 122147 81479 122175
rect 81507 122147 81541 122175
rect 81569 122147 81603 122175
rect 81631 122147 81679 122175
rect 81369 122113 81679 122147
rect 81369 122085 81417 122113
rect 81445 122085 81479 122113
rect 81507 122085 81541 122113
rect 81569 122085 81603 122113
rect 81631 122085 81679 122113
rect 81369 122051 81679 122085
rect 81369 122023 81417 122051
rect 81445 122023 81479 122051
rect 81507 122023 81541 122051
rect 81569 122023 81603 122051
rect 81631 122023 81679 122051
rect 81369 121989 81679 122023
rect 81369 121961 81417 121989
rect 81445 121961 81479 121989
rect 81507 121961 81541 121989
rect 81569 121961 81603 121989
rect 81631 121961 81679 121989
rect 81369 113175 81679 121961
rect 81369 113147 81417 113175
rect 81445 113147 81479 113175
rect 81507 113147 81541 113175
rect 81569 113147 81603 113175
rect 81631 113147 81679 113175
rect 81369 113113 81679 113147
rect 81369 113085 81417 113113
rect 81445 113085 81479 113113
rect 81507 113085 81541 113113
rect 81569 113085 81603 113113
rect 81631 113085 81679 113113
rect 81369 113051 81679 113085
rect 81369 113023 81417 113051
rect 81445 113023 81479 113051
rect 81507 113023 81541 113051
rect 81569 113023 81603 113051
rect 81631 113023 81679 113051
rect 81369 112989 81679 113023
rect 81369 112961 81417 112989
rect 81445 112961 81479 112989
rect 81507 112961 81541 112989
rect 81569 112961 81603 112989
rect 81631 112961 81679 112989
rect 81369 104175 81679 112961
rect 81369 104147 81417 104175
rect 81445 104147 81479 104175
rect 81507 104147 81541 104175
rect 81569 104147 81603 104175
rect 81631 104147 81679 104175
rect 81369 104113 81679 104147
rect 81369 104085 81417 104113
rect 81445 104085 81479 104113
rect 81507 104085 81541 104113
rect 81569 104085 81603 104113
rect 81631 104085 81679 104113
rect 81369 104051 81679 104085
rect 81369 104023 81417 104051
rect 81445 104023 81479 104051
rect 81507 104023 81541 104051
rect 81569 104023 81603 104051
rect 81631 104023 81679 104051
rect 81369 103989 81679 104023
rect 81369 103961 81417 103989
rect 81445 103961 81479 103989
rect 81507 103961 81541 103989
rect 81569 103961 81603 103989
rect 81631 103961 81679 103989
rect 81369 95175 81679 103961
rect 94869 128175 95179 136961
rect 94869 128147 94917 128175
rect 94945 128147 94979 128175
rect 95007 128147 95041 128175
rect 95069 128147 95103 128175
rect 95131 128147 95179 128175
rect 94869 128113 95179 128147
rect 94869 128085 94917 128113
rect 94945 128085 94979 128113
rect 95007 128085 95041 128113
rect 95069 128085 95103 128113
rect 95131 128085 95179 128113
rect 94869 128051 95179 128085
rect 94869 128023 94917 128051
rect 94945 128023 94979 128051
rect 95007 128023 95041 128051
rect 95069 128023 95103 128051
rect 95131 128023 95179 128051
rect 94869 127989 95179 128023
rect 94869 127961 94917 127989
rect 94945 127961 94979 127989
rect 95007 127961 95041 127989
rect 95069 127961 95103 127989
rect 95131 127961 95179 127989
rect 94869 119175 95179 127961
rect 94869 119147 94917 119175
rect 94945 119147 94979 119175
rect 95007 119147 95041 119175
rect 95069 119147 95103 119175
rect 95131 119147 95179 119175
rect 94869 119113 95179 119147
rect 94869 119085 94917 119113
rect 94945 119085 94979 119113
rect 95007 119085 95041 119113
rect 95069 119085 95103 119113
rect 95131 119085 95179 119113
rect 94869 119051 95179 119085
rect 94869 119023 94917 119051
rect 94945 119023 94979 119051
rect 95007 119023 95041 119051
rect 95069 119023 95103 119051
rect 95131 119023 95179 119051
rect 94869 118989 95179 119023
rect 94869 118961 94917 118989
rect 94945 118961 94979 118989
rect 95007 118961 95041 118989
rect 95069 118961 95103 118989
rect 95131 118961 95179 118989
rect 94869 110175 95179 118961
rect 94869 110147 94917 110175
rect 94945 110147 94979 110175
rect 95007 110147 95041 110175
rect 95069 110147 95103 110175
rect 95131 110147 95179 110175
rect 94869 110113 95179 110147
rect 94869 110085 94917 110113
rect 94945 110085 94979 110113
rect 95007 110085 95041 110113
rect 95069 110085 95103 110113
rect 95131 110085 95179 110113
rect 94869 110051 95179 110085
rect 94869 110023 94917 110051
rect 94945 110023 94979 110051
rect 95007 110023 95041 110051
rect 95069 110023 95103 110051
rect 95131 110023 95179 110051
rect 94869 109989 95179 110023
rect 94869 109961 94917 109989
rect 94945 109961 94979 109989
rect 95007 109961 95041 109989
rect 95069 109961 95103 109989
rect 95131 109961 95179 109989
rect 93024 101175 93184 101192
rect 93024 101147 93059 101175
rect 93087 101147 93121 101175
rect 93149 101147 93184 101175
rect 93024 101113 93184 101147
rect 93024 101085 93059 101113
rect 93087 101085 93121 101113
rect 93149 101085 93184 101113
rect 93024 101051 93184 101085
rect 93024 101023 93059 101051
rect 93087 101023 93121 101051
rect 93149 101023 93184 101051
rect 93024 100989 93184 101023
rect 93024 100961 93059 100989
rect 93087 100961 93121 100989
rect 93149 100961 93184 100989
rect 93024 100944 93184 100961
rect 94869 101175 95179 109961
rect 94869 101147 94917 101175
rect 94945 101147 94979 101175
rect 95007 101147 95041 101175
rect 95069 101147 95103 101175
rect 95131 101147 95179 101175
rect 94869 101113 95179 101147
rect 94869 101085 94917 101113
rect 94945 101085 94979 101113
rect 95007 101085 95041 101113
rect 95069 101085 95103 101113
rect 95131 101085 95179 101113
rect 94869 101051 95179 101085
rect 94869 101023 94917 101051
rect 94945 101023 94979 101051
rect 95007 101023 95041 101051
rect 95069 101023 95103 101051
rect 95131 101023 95179 101051
rect 94869 100989 95179 101023
rect 94869 100961 94917 100989
rect 94945 100961 94979 100989
rect 95007 100961 95041 100989
rect 95069 100961 95103 100989
rect 95131 100961 95179 100989
rect 81369 95147 81417 95175
rect 81445 95147 81479 95175
rect 81507 95147 81541 95175
rect 81569 95147 81603 95175
rect 81631 95147 81679 95175
rect 81369 95113 81679 95147
rect 81369 95085 81417 95113
rect 81445 95085 81479 95113
rect 81507 95085 81541 95113
rect 81569 95085 81603 95113
rect 81631 95085 81679 95113
rect 81369 95051 81679 95085
rect 81369 95023 81417 95051
rect 81445 95023 81479 95051
rect 81507 95023 81541 95051
rect 81569 95023 81603 95051
rect 81631 95023 81679 95051
rect 81369 94989 81679 95023
rect 81369 94961 81417 94989
rect 81445 94961 81479 94989
rect 81507 94961 81541 94989
rect 81569 94961 81603 94989
rect 81631 94961 81679 94989
rect 81369 86175 81679 94961
rect 85344 95175 85504 95192
rect 85344 95147 85379 95175
rect 85407 95147 85441 95175
rect 85469 95147 85504 95175
rect 85344 95113 85504 95147
rect 85344 95085 85379 95113
rect 85407 95085 85441 95113
rect 85469 95085 85504 95113
rect 85344 95051 85504 95085
rect 85344 95023 85379 95051
rect 85407 95023 85441 95051
rect 85469 95023 85504 95051
rect 85344 94989 85504 95023
rect 85344 94961 85379 94989
rect 85407 94961 85441 94989
rect 85469 94961 85504 94989
rect 85344 94944 85504 94961
rect 93024 92175 93184 92192
rect 93024 92147 93059 92175
rect 93087 92147 93121 92175
rect 93149 92147 93184 92175
rect 93024 92113 93184 92147
rect 93024 92085 93059 92113
rect 93087 92085 93121 92113
rect 93149 92085 93184 92113
rect 93024 92051 93184 92085
rect 93024 92023 93059 92051
rect 93087 92023 93121 92051
rect 93149 92023 93184 92051
rect 93024 91989 93184 92023
rect 93024 91961 93059 91989
rect 93087 91961 93121 91989
rect 93149 91961 93184 91989
rect 93024 91944 93184 91961
rect 94869 92175 95179 100961
rect 94869 92147 94917 92175
rect 94945 92147 94979 92175
rect 95007 92147 95041 92175
rect 95069 92147 95103 92175
rect 95131 92147 95179 92175
rect 94869 92113 95179 92147
rect 94869 92085 94917 92113
rect 94945 92085 94979 92113
rect 95007 92085 95041 92113
rect 95069 92085 95103 92113
rect 95131 92085 95179 92113
rect 94869 92051 95179 92085
rect 94869 92023 94917 92051
rect 94945 92023 94979 92051
rect 95007 92023 95041 92051
rect 95069 92023 95103 92051
rect 95131 92023 95179 92051
rect 94869 91989 95179 92023
rect 94869 91961 94917 91989
rect 94945 91961 94979 91989
rect 95007 91961 95041 91989
rect 95069 91961 95103 91989
rect 95131 91961 95179 91989
rect 81369 86147 81417 86175
rect 81445 86147 81479 86175
rect 81507 86147 81541 86175
rect 81569 86147 81603 86175
rect 81631 86147 81679 86175
rect 81369 86113 81679 86147
rect 81369 86085 81417 86113
rect 81445 86085 81479 86113
rect 81507 86085 81541 86113
rect 81569 86085 81603 86113
rect 81631 86085 81679 86113
rect 81369 86051 81679 86085
rect 81369 86023 81417 86051
rect 81445 86023 81479 86051
rect 81507 86023 81541 86051
rect 81569 86023 81603 86051
rect 81631 86023 81679 86051
rect 81369 85989 81679 86023
rect 81369 85961 81417 85989
rect 81445 85961 81479 85989
rect 81507 85961 81541 85989
rect 81569 85961 81603 85989
rect 81631 85961 81679 85989
rect 81369 77175 81679 85961
rect 85344 86175 85504 86192
rect 85344 86147 85379 86175
rect 85407 86147 85441 86175
rect 85469 86147 85504 86175
rect 85344 86113 85504 86147
rect 85344 86085 85379 86113
rect 85407 86085 85441 86113
rect 85469 86085 85504 86113
rect 85344 86051 85504 86085
rect 85344 86023 85379 86051
rect 85407 86023 85441 86051
rect 85469 86023 85504 86051
rect 85344 85989 85504 86023
rect 85344 85961 85379 85989
rect 85407 85961 85441 85989
rect 85469 85961 85504 85989
rect 85344 85944 85504 85961
rect 93024 83175 93184 83192
rect 93024 83147 93059 83175
rect 93087 83147 93121 83175
rect 93149 83147 93184 83175
rect 93024 83113 93184 83147
rect 93024 83085 93059 83113
rect 93087 83085 93121 83113
rect 93149 83085 93184 83113
rect 93024 83051 93184 83085
rect 93024 83023 93059 83051
rect 93087 83023 93121 83051
rect 93149 83023 93184 83051
rect 93024 82989 93184 83023
rect 93024 82961 93059 82989
rect 93087 82961 93121 82989
rect 93149 82961 93184 82989
rect 93024 82944 93184 82961
rect 94869 83175 95179 91961
rect 94869 83147 94917 83175
rect 94945 83147 94979 83175
rect 95007 83147 95041 83175
rect 95069 83147 95103 83175
rect 95131 83147 95179 83175
rect 94869 83113 95179 83147
rect 94869 83085 94917 83113
rect 94945 83085 94979 83113
rect 95007 83085 95041 83113
rect 95069 83085 95103 83113
rect 95131 83085 95179 83113
rect 94869 83051 95179 83085
rect 94869 83023 94917 83051
rect 94945 83023 94979 83051
rect 95007 83023 95041 83051
rect 95069 83023 95103 83051
rect 95131 83023 95179 83051
rect 94869 82989 95179 83023
rect 94869 82961 94917 82989
rect 94945 82961 94979 82989
rect 95007 82961 95041 82989
rect 95069 82961 95103 82989
rect 95131 82961 95179 82989
rect 81369 77147 81417 77175
rect 81445 77147 81479 77175
rect 81507 77147 81541 77175
rect 81569 77147 81603 77175
rect 81631 77147 81679 77175
rect 81369 77113 81679 77147
rect 81369 77085 81417 77113
rect 81445 77085 81479 77113
rect 81507 77085 81541 77113
rect 81569 77085 81603 77113
rect 81631 77085 81679 77113
rect 81369 77051 81679 77085
rect 81369 77023 81417 77051
rect 81445 77023 81479 77051
rect 81507 77023 81541 77051
rect 81569 77023 81603 77051
rect 81631 77023 81679 77051
rect 81369 76989 81679 77023
rect 81369 76961 81417 76989
rect 81445 76961 81479 76989
rect 81507 76961 81541 76989
rect 81569 76961 81603 76989
rect 81631 76961 81679 76989
rect 81369 68175 81679 76961
rect 85344 77175 85504 77192
rect 85344 77147 85379 77175
rect 85407 77147 85441 77175
rect 85469 77147 85504 77175
rect 85344 77113 85504 77147
rect 85344 77085 85379 77113
rect 85407 77085 85441 77113
rect 85469 77085 85504 77113
rect 85344 77051 85504 77085
rect 85344 77023 85379 77051
rect 85407 77023 85441 77051
rect 85469 77023 85504 77051
rect 85344 76989 85504 77023
rect 85344 76961 85379 76989
rect 85407 76961 85441 76989
rect 85469 76961 85504 76989
rect 85344 76944 85504 76961
rect 81369 68147 81417 68175
rect 81445 68147 81479 68175
rect 81507 68147 81541 68175
rect 81569 68147 81603 68175
rect 81631 68147 81679 68175
rect 81369 68113 81679 68147
rect 81369 68085 81417 68113
rect 81445 68085 81479 68113
rect 81507 68085 81541 68113
rect 81569 68085 81603 68113
rect 81631 68085 81679 68113
rect 81369 68051 81679 68085
rect 81369 68023 81417 68051
rect 81445 68023 81479 68051
rect 81507 68023 81541 68051
rect 81569 68023 81603 68051
rect 81631 68023 81679 68051
rect 81369 67989 81679 68023
rect 81369 67961 81417 67989
rect 81445 67961 81479 67989
rect 81507 67961 81541 67989
rect 81569 67961 81603 67989
rect 81631 67961 81679 67989
rect 81369 59175 81679 67961
rect 81369 59147 81417 59175
rect 81445 59147 81479 59175
rect 81507 59147 81541 59175
rect 81569 59147 81603 59175
rect 81631 59147 81679 59175
rect 81369 59113 81679 59147
rect 81369 59085 81417 59113
rect 81445 59085 81479 59113
rect 81507 59085 81541 59113
rect 81569 59085 81603 59113
rect 81631 59085 81679 59113
rect 81369 59051 81679 59085
rect 81369 59023 81417 59051
rect 81445 59023 81479 59051
rect 81507 59023 81541 59051
rect 81569 59023 81603 59051
rect 81631 59023 81679 59051
rect 81369 58989 81679 59023
rect 81369 58961 81417 58989
rect 81445 58961 81479 58989
rect 81507 58961 81541 58989
rect 81569 58961 81603 58989
rect 81631 58961 81679 58989
rect 81369 50175 81679 58961
rect 81369 50147 81417 50175
rect 81445 50147 81479 50175
rect 81507 50147 81541 50175
rect 81569 50147 81603 50175
rect 81631 50147 81679 50175
rect 81369 50113 81679 50147
rect 81369 50085 81417 50113
rect 81445 50085 81479 50113
rect 81507 50085 81541 50113
rect 81569 50085 81603 50113
rect 81631 50085 81679 50113
rect 81369 50051 81679 50085
rect 81369 50023 81417 50051
rect 81445 50023 81479 50051
rect 81507 50023 81541 50051
rect 81569 50023 81603 50051
rect 81631 50023 81679 50051
rect 81369 49989 81679 50023
rect 81369 49961 81417 49989
rect 81445 49961 81479 49989
rect 81507 49961 81541 49989
rect 81569 49961 81603 49989
rect 81631 49961 81679 49989
rect 81369 41175 81679 49961
rect 81369 41147 81417 41175
rect 81445 41147 81479 41175
rect 81507 41147 81541 41175
rect 81569 41147 81603 41175
rect 81631 41147 81679 41175
rect 81369 41113 81679 41147
rect 81369 41085 81417 41113
rect 81445 41085 81479 41113
rect 81507 41085 81541 41113
rect 81569 41085 81603 41113
rect 81631 41085 81679 41113
rect 81369 41051 81679 41085
rect 81369 41023 81417 41051
rect 81445 41023 81479 41051
rect 81507 41023 81541 41051
rect 81569 41023 81603 41051
rect 81631 41023 81679 41051
rect 81369 40989 81679 41023
rect 81369 40961 81417 40989
rect 81445 40961 81479 40989
rect 81507 40961 81541 40989
rect 81569 40961 81603 40989
rect 81631 40961 81679 40989
rect 81369 32175 81679 40961
rect 81369 32147 81417 32175
rect 81445 32147 81479 32175
rect 81507 32147 81541 32175
rect 81569 32147 81603 32175
rect 81631 32147 81679 32175
rect 81369 32113 81679 32147
rect 81369 32085 81417 32113
rect 81445 32085 81479 32113
rect 81507 32085 81541 32113
rect 81569 32085 81603 32113
rect 81631 32085 81679 32113
rect 81369 32051 81679 32085
rect 81369 32023 81417 32051
rect 81445 32023 81479 32051
rect 81507 32023 81541 32051
rect 81569 32023 81603 32051
rect 81631 32023 81679 32051
rect 81369 31989 81679 32023
rect 81369 31961 81417 31989
rect 81445 31961 81479 31989
rect 81507 31961 81541 31989
rect 81569 31961 81603 31989
rect 81631 31961 81679 31989
rect 81369 23175 81679 31961
rect 81369 23147 81417 23175
rect 81445 23147 81479 23175
rect 81507 23147 81541 23175
rect 81569 23147 81603 23175
rect 81631 23147 81679 23175
rect 81369 23113 81679 23147
rect 81369 23085 81417 23113
rect 81445 23085 81479 23113
rect 81507 23085 81541 23113
rect 81569 23085 81603 23113
rect 81631 23085 81679 23113
rect 81369 23051 81679 23085
rect 81369 23023 81417 23051
rect 81445 23023 81479 23051
rect 81507 23023 81541 23051
rect 81569 23023 81603 23051
rect 81631 23023 81679 23051
rect 81369 22989 81679 23023
rect 81369 22961 81417 22989
rect 81445 22961 81479 22989
rect 81507 22961 81541 22989
rect 81569 22961 81603 22989
rect 81631 22961 81679 22989
rect 81369 14175 81679 22961
rect 81369 14147 81417 14175
rect 81445 14147 81479 14175
rect 81507 14147 81541 14175
rect 81569 14147 81603 14175
rect 81631 14147 81679 14175
rect 81369 14113 81679 14147
rect 81369 14085 81417 14113
rect 81445 14085 81479 14113
rect 81507 14085 81541 14113
rect 81569 14085 81603 14113
rect 81631 14085 81679 14113
rect 81369 14051 81679 14085
rect 81369 14023 81417 14051
rect 81445 14023 81479 14051
rect 81507 14023 81541 14051
rect 81569 14023 81603 14051
rect 81631 14023 81679 14051
rect 81369 13989 81679 14023
rect 81369 13961 81417 13989
rect 81445 13961 81479 13989
rect 81507 13961 81541 13989
rect 81569 13961 81603 13989
rect 81631 13961 81679 13989
rect 81369 5175 81679 13961
rect 81369 5147 81417 5175
rect 81445 5147 81479 5175
rect 81507 5147 81541 5175
rect 81569 5147 81603 5175
rect 81631 5147 81679 5175
rect 81369 5113 81679 5147
rect 81369 5085 81417 5113
rect 81445 5085 81479 5113
rect 81507 5085 81541 5113
rect 81569 5085 81603 5113
rect 81631 5085 81679 5113
rect 81369 5051 81679 5085
rect 81369 5023 81417 5051
rect 81445 5023 81479 5051
rect 81507 5023 81541 5051
rect 81569 5023 81603 5051
rect 81631 5023 81679 5051
rect 81369 4989 81679 5023
rect 81369 4961 81417 4989
rect 81445 4961 81479 4989
rect 81507 4961 81541 4989
rect 81569 4961 81603 4989
rect 81631 4961 81679 4989
rect 81369 -560 81679 4961
rect 81369 -588 81417 -560
rect 81445 -588 81479 -560
rect 81507 -588 81541 -560
rect 81569 -588 81603 -560
rect 81631 -588 81679 -560
rect 81369 -622 81679 -588
rect 81369 -650 81417 -622
rect 81445 -650 81479 -622
rect 81507 -650 81541 -622
rect 81569 -650 81603 -622
rect 81631 -650 81679 -622
rect 81369 -684 81679 -650
rect 81369 -712 81417 -684
rect 81445 -712 81479 -684
rect 81507 -712 81541 -684
rect 81569 -712 81603 -684
rect 81631 -712 81679 -684
rect 81369 -746 81679 -712
rect 81369 -774 81417 -746
rect 81445 -774 81479 -746
rect 81507 -774 81541 -746
rect 81569 -774 81603 -746
rect 81631 -774 81679 -746
rect 81369 -822 81679 -774
rect 94869 74175 95179 82961
rect 94869 74147 94917 74175
rect 94945 74147 94979 74175
rect 95007 74147 95041 74175
rect 95069 74147 95103 74175
rect 95131 74147 95179 74175
rect 94869 74113 95179 74147
rect 94869 74085 94917 74113
rect 94945 74085 94979 74113
rect 95007 74085 95041 74113
rect 95069 74085 95103 74113
rect 95131 74085 95179 74113
rect 94869 74051 95179 74085
rect 94869 74023 94917 74051
rect 94945 74023 94979 74051
rect 95007 74023 95041 74051
rect 95069 74023 95103 74051
rect 95131 74023 95179 74051
rect 94869 73989 95179 74023
rect 94869 73961 94917 73989
rect 94945 73961 94979 73989
rect 95007 73961 95041 73989
rect 95069 73961 95103 73989
rect 95131 73961 95179 73989
rect 94869 65175 95179 73961
rect 94869 65147 94917 65175
rect 94945 65147 94979 65175
rect 95007 65147 95041 65175
rect 95069 65147 95103 65175
rect 95131 65147 95179 65175
rect 94869 65113 95179 65147
rect 94869 65085 94917 65113
rect 94945 65085 94979 65113
rect 95007 65085 95041 65113
rect 95069 65085 95103 65113
rect 95131 65085 95179 65113
rect 94869 65051 95179 65085
rect 94869 65023 94917 65051
rect 94945 65023 94979 65051
rect 95007 65023 95041 65051
rect 95069 65023 95103 65051
rect 95131 65023 95179 65051
rect 94869 64989 95179 65023
rect 94869 64961 94917 64989
rect 94945 64961 94979 64989
rect 95007 64961 95041 64989
rect 95069 64961 95103 64989
rect 95131 64961 95179 64989
rect 94869 56175 95179 64961
rect 94869 56147 94917 56175
rect 94945 56147 94979 56175
rect 95007 56147 95041 56175
rect 95069 56147 95103 56175
rect 95131 56147 95179 56175
rect 94869 56113 95179 56147
rect 94869 56085 94917 56113
rect 94945 56085 94979 56113
rect 95007 56085 95041 56113
rect 95069 56085 95103 56113
rect 95131 56085 95179 56113
rect 94869 56051 95179 56085
rect 94869 56023 94917 56051
rect 94945 56023 94979 56051
rect 95007 56023 95041 56051
rect 95069 56023 95103 56051
rect 95131 56023 95179 56051
rect 94869 55989 95179 56023
rect 94869 55961 94917 55989
rect 94945 55961 94979 55989
rect 95007 55961 95041 55989
rect 95069 55961 95103 55989
rect 95131 55961 95179 55989
rect 94869 47175 95179 55961
rect 94869 47147 94917 47175
rect 94945 47147 94979 47175
rect 95007 47147 95041 47175
rect 95069 47147 95103 47175
rect 95131 47147 95179 47175
rect 94869 47113 95179 47147
rect 94869 47085 94917 47113
rect 94945 47085 94979 47113
rect 95007 47085 95041 47113
rect 95069 47085 95103 47113
rect 95131 47085 95179 47113
rect 94869 47051 95179 47085
rect 94869 47023 94917 47051
rect 94945 47023 94979 47051
rect 95007 47023 95041 47051
rect 95069 47023 95103 47051
rect 95131 47023 95179 47051
rect 94869 46989 95179 47023
rect 94869 46961 94917 46989
rect 94945 46961 94979 46989
rect 95007 46961 95041 46989
rect 95069 46961 95103 46989
rect 95131 46961 95179 46989
rect 94869 38175 95179 46961
rect 94869 38147 94917 38175
rect 94945 38147 94979 38175
rect 95007 38147 95041 38175
rect 95069 38147 95103 38175
rect 95131 38147 95179 38175
rect 94869 38113 95179 38147
rect 94869 38085 94917 38113
rect 94945 38085 94979 38113
rect 95007 38085 95041 38113
rect 95069 38085 95103 38113
rect 95131 38085 95179 38113
rect 94869 38051 95179 38085
rect 94869 38023 94917 38051
rect 94945 38023 94979 38051
rect 95007 38023 95041 38051
rect 95069 38023 95103 38051
rect 95131 38023 95179 38051
rect 94869 37989 95179 38023
rect 94869 37961 94917 37989
rect 94945 37961 94979 37989
rect 95007 37961 95041 37989
rect 95069 37961 95103 37989
rect 95131 37961 95179 37989
rect 94869 29175 95179 37961
rect 94869 29147 94917 29175
rect 94945 29147 94979 29175
rect 95007 29147 95041 29175
rect 95069 29147 95103 29175
rect 95131 29147 95179 29175
rect 94869 29113 95179 29147
rect 94869 29085 94917 29113
rect 94945 29085 94979 29113
rect 95007 29085 95041 29113
rect 95069 29085 95103 29113
rect 95131 29085 95179 29113
rect 94869 29051 95179 29085
rect 94869 29023 94917 29051
rect 94945 29023 94979 29051
rect 95007 29023 95041 29051
rect 95069 29023 95103 29051
rect 95131 29023 95179 29051
rect 94869 28989 95179 29023
rect 94869 28961 94917 28989
rect 94945 28961 94979 28989
rect 95007 28961 95041 28989
rect 95069 28961 95103 28989
rect 95131 28961 95179 28989
rect 94869 20175 95179 28961
rect 94869 20147 94917 20175
rect 94945 20147 94979 20175
rect 95007 20147 95041 20175
rect 95069 20147 95103 20175
rect 95131 20147 95179 20175
rect 94869 20113 95179 20147
rect 94869 20085 94917 20113
rect 94945 20085 94979 20113
rect 95007 20085 95041 20113
rect 95069 20085 95103 20113
rect 95131 20085 95179 20113
rect 94869 20051 95179 20085
rect 94869 20023 94917 20051
rect 94945 20023 94979 20051
rect 95007 20023 95041 20051
rect 95069 20023 95103 20051
rect 95131 20023 95179 20051
rect 94869 19989 95179 20023
rect 94869 19961 94917 19989
rect 94945 19961 94979 19989
rect 95007 19961 95041 19989
rect 95069 19961 95103 19989
rect 95131 19961 95179 19989
rect 94869 11175 95179 19961
rect 94869 11147 94917 11175
rect 94945 11147 94979 11175
rect 95007 11147 95041 11175
rect 95069 11147 95103 11175
rect 95131 11147 95179 11175
rect 94869 11113 95179 11147
rect 94869 11085 94917 11113
rect 94945 11085 94979 11113
rect 95007 11085 95041 11113
rect 95069 11085 95103 11113
rect 95131 11085 95179 11113
rect 94869 11051 95179 11085
rect 94869 11023 94917 11051
rect 94945 11023 94979 11051
rect 95007 11023 95041 11051
rect 95069 11023 95103 11051
rect 95131 11023 95179 11051
rect 94869 10989 95179 11023
rect 94869 10961 94917 10989
rect 94945 10961 94979 10989
rect 95007 10961 95041 10989
rect 95069 10961 95103 10989
rect 95131 10961 95179 10989
rect 94869 2175 95179 10961
rect 94869 2147 94917 2175
rect 94945 2147 94979 2175
rect 95007 2147 95041 2175
rect 95069 2147 95103 2175
rect 95131 2147 95179 2175
rect 94869 2113 95179 2147
rect 94869 2085 94917 2113
rect 94945 2085 94979 2113
rect 95007 2085 95041 2113
rect 95069 2085 95103 2113
rect 95131 2085 95179 2113
rect 94869 2051 95179 2085
rect 94869 2023 94917 2051
rect 94945 2023 94979 2051
rect 95007 2023 95041 2051
rect 95069 2023 95103 2051
rect 95131 2023 95179 2051
rect 94869 1989 95179 2023
rect 94869 1961 94917 1989
rect 94945 1961 94979 1989
rect 95007 1961 95041 1989
rect 95069 1961 95103 1989
rect 95131 1961 95179 1989
rect 94869 -80 95179 1961
rect 94869 -108 94917 -80
rect 94945 -108 94979 -80
rect 95007 -108 95041 -80
rect 95069 -108 95103 -80
rect 95131 -108 95179 -80
rect 94869 -142 95179 -108
rect 94869 -170 94917 -142
rect 94945 -170 94979 -142
rect 95007 -170 95041 -142
rect 95069 -170 95103 -142
rect 95131 -170 95179 -142
rect 94869 -204 95179 -170
rect 94869 -232 94917 -204
rect 94945 -232 94979 -204
rect 95007 -232 95041 -204
rect 95069 -232 95103 -204
rect 95131 -232 95179 -204
rect 94869 -266 95179 -232
rect 94869 -294 94917 -266
rect 94945 -294 94979 -266
rect 95007 -294 95041 -266
rect 95069 -294 95103 -266
rect 95131 -294 95179 -266
rect 94869 -822 95179 -294
rect 96729 299086 97039 299134
rect 96729 299058 96777 299086
rect 96805 299058 96839 299086
rect 96867 299058 96901 299086
rect 96929 299058 96963 299086
rect 96991 299058 97039 299086
rect 96729 299024 97039 299058
rect 96729 298996 96777 299024
rect 96805 298996 96839 299024
rect 96867 298996 96901 299024
rect 96929 298996 96963 299024
rect 96991 298996 97039 299024
rect 96729 298962 97039 298996
rect 96729 298934 96777 298962
rect 96805 298934 96839 298962
rect 96867 298934 96901 298962
rect 96929 298934 96963 298962
rect 96991 298934 97039 298962
rect 96729 298900 97039 298934
rect 96729 298872 96777 298900
rect 96805 298872 96839 298900
rect 96867 298872 96901 298900
rect 96929 298872 96963 298900
rect 96991 298872 97039 298900
rect 96729 293175 97039 298872
rect 96729 293147 96777 293175
rect 96805 293147 96839 293175
rect 96867 293147 96901 293175
rect 96929 293147 96963 293175
rect 96991 293147 97039 293175
rect 96729 293113 97039 293147
rect 96729 293085 96777 293113
rect 96805 293085 96839 293113
rect 96867 293085 96901 293113
rect 96929 293085 96963 293113
rect 96991 293085 97039 293113
rect 96729 293051 97039 293085
rect 96729 293023 96777 293051
rect 96805 293023 96839 293051
rect 96867 293023 96901 293051
rect 96929 293023 96963 293051
rect 96991 293023 97039 293051
rect 96729 292989 97039 293023
rect 96729 292961 96777 292989
rect 96805 292961 96839 292989
rect 96867 292961 96901 292989
rect 96929 292961 96963 292989
rect 96991 292961 97039 292989
rect 96729 284175 97039 292961
rect 96729 284147 96777 284175
rect 96805 284147 96839 284175
rect 96867 284147 96901 284175
rect 96929 284147 96963 284175
rect 96991 284147 97039 284175
rect 96729 284113 97039 284147
rect 96729 284085 96777 284113
rect 96805 284085 96839 284113
rect 96867 284085 96901 284113
rect 96929 284085 96963 284113
rect 96991 284085 97039 284113
rect 96729 284051 97039 284085
rect 96729 284023 96777 284051
rect 96805 284023 96839 284051
rect 96867 284023 96901 284051
rect 96929 284023 96963 284051
rect 96991 284023 97039 284051
rect 96729 283989 97039 284023
rect 96729 283961 96777 283989
rect 96805 283961 96839 283989
rect 96867 283961 96901 283989
rect 96929 283961 96963 283989
rect 96991 283961 97039 283989
rect 96729 275175 97039 283961
rect 96729 275147 96777 275175
rect 96805 275147 96839 275175
rect 96867 275147 96901 275175
rect 96929 275147 96963 275175
rect 96991 275147 97039 275175
rect 96729 275113 97039 275147
rect 96729 275085 96777 275113
rect 96805 275085 96839 275113
rect 96867 275085 96901 275113
rect 96929 275085 96963 275113
rect 96991 275085 97039 275113
rect 96729 275051 97039 275085
rect 96729 275023 96777 275051
rect 96805 275023 96839 275051
rect 96867 275023 96901 275051
rect 96929 275023 96963 275051
rect 96991 275023 97039 275051
rect 96729 274989 97039 275023
rect 96729 274961 96777 274989
rect 96805 274961 96839 274989
rect 96867 274961 96901 274989
rect 96929 274961 96963 274989
rect 96991 274961 97039 274989
rect 96729 266175 97039 274961
rect 110229 298606 110539 299134
rect 110229 298578 110277 298606
rect 110305 298578 110339 298606
rect 110367 298578 110401 298606
rect 110429 298578 110463 298606
rect 110491 298578 110539 298606
rect 110229 298544 110539 298578
rect 110229 298516 110277 298544
rect 110305 298516 110339 298544
rect 110367 298516 110401 298544
rect 110429 298516 110463 298544
rect 110491 298516 110539 298544
rect 110229 298482 110539 298516
rect 110229 298454 110277 298482
rect 110305 298454 110339 298482
rect 110367 298454 110401 298482
rect 110429 298454 110463 298482
rect 110491 298454 110539 298482
rect 110229 298420 110539 298454
rect 110229 298392 110277 298420
rect 110305 298392 110339 298420
rect 110367 298392 110401 298420
rect 110429 298392 110463 298420
rect 110491 298392 110539 298420
rect 110229 290175 110539 298392
rect 110229 290147 110277 290175
rect 110305 290147 110339 290175
rect 110367 290147 110401 290175
rect 110429 290147 110463 290175
rect 110491 290147 110539 290175
rect 110229 290113 110539 290147
rect 110229 290085 110277 290113
rect 110305 290085 110339 290113
rect 110367 290085 110401 290113
rect 110429 290085 110463 290113
rect 110491 290085 110539 290113
rect 110229 290051 110539 290085
rect 110229 290023 110277 290051
rect 110305 290023 110339 290051
rect 110367 290023 110401 290051
rect 110429 290023 110463 290051
rect 110491 290023 110539 290051
rect 110229 289989 110539 290023
rect 110229 289961 110277 289989
rect 110305 289961 110339 289989
rect 110367 289961 110401 289989
rect 110429 289961 110463 289989
rect 110491 289961 110539 289989
rect 110229 281175 110539 289961
rect 110229 281147 110277 281175
rect 110305 281147 110339 281175
rect 110367 281147 110401 281175
rect 110429 281147 110463 281175
rect 110491 281147 110539 281175
rect 110229 281113 110539 281147
rect 110229 281085 110277 281113
rect 110305 281085 110339 281113
rect 110367 281085 110401 281113
rect 110429 281085 110463 281113
rect 110491 281085 110539 281113
rect 110229 281051 110539 281085
rect 110229 281023 110277 281051
rect 110305 281023 110339 281051
rect 110367 281023 110401 281051
rect 110429 281023 110463 281051
rect 110491 281023 110539 281051
rect 110229 280989 110539 281023
rect 110229 280961 110277 280989
rect 110305 280961 110339 280989
rect 110367 280961 110401 280989
rect 110429 280961 110463 280989
rect 110491 280961 110539 280989
rect 110229 272175 110539 280961
rect 110229 272147 110277 272175
rect 110305 272147 110339 272175
rect 110367 272147 110401 272175
rect 110429 272147 110463 272175
rect 110491 272147 110539 272175
rect 110229 272113 110539 272147
rect 110229 272085 110277 272113
rect 110305 272085 110339 272113
rect 110367 272085 110401 272113
rect 110429 272085 110463 272113
rect 110491 272085 110539 272113
rect 110229 272051 110539 272085
rect 110229 272023 110277 272051
rect 110305 272023 110339 272051
rect 110367 272023 110401 272051
rect 110429 272023 110463 272051
rect 110491 272023 110539 272051
rect 110229 271989 110539 272023
rect 110229 271961 110277 271989
rect 110305 271961 110339 271989
rect 110367 271961 110401 271989
rect 110429 271961 110463 271989
rect 110491 271961 110539 271989
rect 110229 268935 110539 271961
rect 112089 299086 112399 299134
rect 112089 299058 112137 299086
rect 112165 299058 112199 299086
rect 112227 299058 112261 299086
rect 112289 299058 112323 299086
rect 112351 299058 112399 299086
rect 112089 299024 112399 299058
rect 112089 298996 112137 299024
rect 112165 298996 112199 299024
rect 112227 298996 112261 299024
rect 112289 298996 112323 299024
rect 112351 298996 112399 299024
rect 112089 298962 112399 298996
rect 112089 298934 112137 298962
rect 112165 298934 112199 298962
rect 112227 298934 112261 298962
rect 112289 298934 112323 298962
rect 112351 298934 112399 298962
rect 112089 298900 112399 298934
rect 112089 298872 112137 298900
rect 112165 298872 112199 298900
rect 112227 298872 112261 298900
rect 112289 298872 112323 298900
rect 112351 298872 112399 298900
rect 112089 293175 112399 298872
rect 112089 293147 112137 293175
rect 112165 293147 112199 293175
rect 112227 293147 112261 293175
rect 112289 293147 112323 293175
rect 112351 293147 112399 293175
rect 112089 293113 112399 293147
rect 112089 293085 112137 293113
rect 112165 293085 112199 293113
rect 112227 293085 112261 293113
rect 112289 293085 112323 293113
rect 112351 293085 112399 293113
rect 112089 293051 112399 293085
rect 112089 293023 112137 293051
rect 112165 293023 112199 293051
rect 112227 293023 112261 293051
rect 112289 293023 112323 293051
rect 112351 293023 112399 293051
rect 112089 292989 112399 293023
rect 112089 292961 112137 292989
rect 112165 292961 112199 292989
rect 112227 292961 112261 292989
rect 112289 292961 112323 292989
rect 112351 292961 112399 292989
rect 112089 284175 112399 292961
rect 112089 284147 112137 284175
rect 112165 284147 112199 284175
rect 112227 284147 112261 284175
rect 112289 284147 112323 284175
rect 112351 284147 112399 284175
rect 112089 284113 112399 284147
rect 112089 284085 112137 284113
rect 112165 284085 112199 284113
rect 112227 284085 112261 284113
rect 112289 284085 112323 284113
rect 112351 284085 112399 284113
rect 112089 284051 112399 284085
rect 112089 284023 112137 284051
rect 112165 284023 112199 284051
rect 112227 284023 112261 284051
rect 112289 284023 112323 284051
rect 112351 284023 112399 284051
rect 112089 283989 112399 284023
rect 112089 283961 112137 283989
rect 112165 283961 112199 283989
rect 112227 283961 112261 283989
rect 112289 283961 112323 283989
rect 112351 283961 112399 283989
rect 112089 275175 112399 283961
rect 112089 275147 112137 275175
rect 112165 275147 112199 275175
rect 112227 275147 112261 275175
rect 112289 275147 112323 275175
rect 112351 275147 112399 275175
rect 112089 275113 112399 275147
rect 112089 275085 112137 275113
rect 112165 275085 112199 275113
rect 112227 275085 112261 275113
rect 112289 275085 112323 275113
rect 112351 275085 112399 275113
rect 112089 275051 112399 275085
rect 112089 275023 112137 275051
rect 112165 275023 112199 275051
rect 112227 275023 112261 275051
rect 112289 275023 112323 275051
rect 112351 275023 112399 275051
rect 112089 274989 112399 275023
rect 112089 274961 112137 274989
rect 112165 274961 112199 274989
rect 112227 274961 112261 274989
rect 112289 274961 112323 274989
rect 112351 274961 112399 274989
rect 112089 268935 112399 274961
rect 125589 298606 125899 299134
rect 125589 298578 125637 298606
rect 125665 298578 125699 298606
rect 125727 298578 125761 298606
rect 125789 298578 125823 298606
rect 125851 298578 125899 298606
rect 125589 298544 125899 298578
rect 125589 298516 125637 298544
rect 125665 298516 125699 298544
rect 125727 298516 125761 298544
rect 125789 298516 125823 298544
rect 125851 298516 125899 298544
rect 125589 298482 125899 298516
rect 125589 298454 125637 298482
rect 125665 298454 125699 298482
rect 125727 298454 125761 298482
rect 125789 298454 125823 298482
rect 125851 298454 125899 298482
rect 125589 298420 125899 298454
rect 125589 298392 125637 298420
rect 125665 298392 125699 298420
rect 125727 298392 125761 298420
rect 125789 298392 125823 298420
rect 125851 298392 125899 298420
rect 125589 290175 125899 298392
rect 125589 290147 125637 290175
rect 125665 290147 125699 290175
rect 125727 290147 125761 290175
rect 125789 290147 125823 290175
rect 125851 290147 125899 290175
rect 125589 290113 125899 290147
rect 125589 290085 125637 290113
rect 125665 290085 125699 290113
rect 125727 290085 125761 290113
rect 125789 290085 125823 290113
rect 125851 290085 125899 290113
rect 125589 290051 125899 290085
rect 125589 290023 125637 290051
rect 125665 290023 125699 290051
rect 125727 290023 125761 290051
rect 125789 290023 125823 290051
rect 125851 290023 125899 290051
rect 125589 289989 125899 290023
rect 125589 289961 125637 289989
rect 125665 289961 125699 289989
rect 125727 289961 125761 289989
rect 125789 289961 125823 289989
rect 125851 289961 125899 289989
rect 125589 281175 125899 289961
rect 125589 281147 125637 281175
rect 125665 281147 125699 281175
rect 125727 281147 125761 281175
rect 125789 281147 125823 281175
rect 125851 281147 125899 281175
rect 125589 281113 125899 281147
rect 125589 281085 125637 281113
rect 125665 281085 125699 281113
rect 125727 281085 125761 281113
rect 125789 281085 125823 281113
rect 125851 281085 125899 281113
rect 125589 281051 125899 281085
rect 125589 281023 125637 281051
rect 125665 281023 125699 281051
rect 125727 281023 125761 281051
rect 125789 281023 125823 281051
rect 125851 281023 125899 281051
rect 125589 280989 125899 281023
rect 125589 280961 125637 280989
rect 125665 280961 125699 280989
rect 125727 280961 125761 280989
rect 125789 280961 125823 280989
rect 125851 280961 125899 280989
rect 125589 272175 125899 280961
rect 125589 272147 125637 272175
rect 125665 272147 125699 272175
rect 125727 272147 125761 272175
rect 125789 272147 125823 272175
rect 125851 272147 125899 272175
rect 125589 272113 125899 272147
rect 125589 272085 125637 272113
rect 125665 272085 125699 272113
rect 125727 272085 125761 272113
rect 125789 272085 125823 272113
rect 125851 272085 125899 272113
rect 125589 272051 125899 272085
rect 125589 272023 125637 272051
rect 125665 272023 125699 272051
rect 125727 272023 125761 272051
rect 125789 272023 125823 272051
rect 125851 272023 125899 272051
rect 125589 271989 125899 272023
rect 125589 271961 125637 271989
rect 125665 271961 125699 271989
rect 125727 271961 125761 271989
rect 125789 271961 125823 271989
rect 125851 271961 125899 271989
rect 125589 268935 125899 271961
rect 127449 299086 127759 299134
rect 127449 299058 127497 299086
rect 127525 299058 127559 299086
rect 127587 299058 127621 299086
rect 127649 299058 127683 299086
rect 127711 299058 127759 299086
rect 127449 299024 127759 299058
rect 127449 298996 127497 299024
rect 127525 298996 127559 299024
rect 127587 298996 127621 299024
rect 127649 298996 127683 299024
rect 127711 298996 127759 299024
rect 127449 298962 127759 298996
rect 127449 298934 127497 298962
rect 127525 298934 127559 298962
rect 127587 298934 127621 298962
rect 127649 298934 127683 298962
rect 127711 298934 127759 298962
rect 127449 298900 127759 298934
rect 127449 298872 127497 298900
rect 127525 298872 127559 298900
rect 127587 298872 127621 298900
rect 127649 298872 127683 298900
rect 127711 298872 127759 298900
rect 127449 293175 127759 298872
rect 127449 293147 127497 293175
rect 127525 293147 127559 293175
rect 127587 293147 127621 293175
rect 127649 293147 127683 293175
rect 127711 293147 127759 293175
rect 127449 293113 127759 293147
rect 127449 293085 127497 293113
rect 127525 293085 127559 293113
rect 127587 293085 127621 293113
rect 127649 293085 127683 293113
rect 127711 293085 127759 293113
rect 127449 293051 127759 293085
rect 127449 293023 127497 293051
rect 127525 293023 127559 293051
rect 127587 293023 127621 293051
rect 127649 293023 127683 293051
rect 127711 293023 127759 293051
rect 127449 292989 127759 293023
rect 127449 292961 127497 292989
rect 127525 292961 127559 292989
rect 127587 292961 127621 292989
rect 127649 292961 127683 292989
rect 127711 292961 127759 292989
rect 127449 284175 127759 292961
rect 127449 284147 127497 284175
rect 127525 284147 127559 284175
rect 127587 284147 127621 284175
rect 127649 284147 127683 284175
rect 127711 284147 127759 284175
rect 127449 284113 127759 284147
rect 127449 284085 127497 284113
rect 127525 284085 127559 284113
rect 127587 284085 127621 284113
rect 127649 284085 127683 284113
rect 127711 284085 127759 284113
rect 127449 284051 127759 284085
rect 127449 284023 127497 284051
rect 127525 284023 127559 284051
rect 127587 284023 127621 284051
rect 127649 284023 127683 284051
rect 127711 284023 127759 284051
rect 127449 283989 127759 284023
rect 127449 283961 127497 283989
rect 127525 283961 127559 283989
rect 127587 283961 127621 283989
rect 127649 283961 127683 283989
rect 127711 283961 127759 283989
rect 127449 275175 127759 283961
rect 127449 275147 127497 275175
rect 127525 275147 127559 275175
rect 127587 275147 127621 275175
rect 127649 275147 127683 275175
rect 127711 275147 127759 275175
rect 127449 275113 127759 275147
rect 127449 275085 127497 275113
rect 127525 275085 127559 275113
rect 127587 275085 127621 275113
rect 127649 275085 127683 275113
rect 127711 275085 127759 275113
rect 127449 275051 127759 275085
rect 127449 275023 127497 275051
rect 127525 275023 127559 275051
rect 127587 275023 127621 275051
rect 127649 275023 127683 275051
rect 127711 275023 127759 275051
rect 127449 274989 127759 275023
rect 127449 274961 127497 274989
rect 127525 274961 127559 274989
rect 127587 274961 127621 274989
rect 127649 274961 127683 274989
rect 127711 274961 127759 274989
rect 127449 268935 127759 274961
rect 140949 298606 141259 299134
rect 140949 298578 140997 298606
rect 141025 298578 141059 298606
rect 141087 298578 141121 298606
rect 141149 298578 141183 298606
rect 141211 298578 141259 298606
rect 140949 298544 141259 298578
rect 140949 298516 140997 298544
rect 141025 298516 141059 298544
rect 141087 298516 141121 298544
rect 141149 298516 141183 298544
rect 141211 298516 141259 298544
rect 140949 298482 141259 298516
rect 140949 298454 140997 298482
rect 141025 298454 141059 298482
rect 141087 298454 141121 298482
rect 141149 298454 141183 298482
rect 141211 298454 141259 298482
rect 140949 298420 141259 298454
rect 140949 298392 140997 298420
rect 141025 298392 141059 298420
rect 141087 298392 141121 298420
rect 141149 298392 141183 298420
rect 141211 298392 141259 298420
rect 140949 290175 141259 298392
rect 140949 290147 140997 290175
rect 141025 290147 141059 290175
rect 141087 290147 141121 290175
rect 141149 290147 141183 290175
rect 141211 290147 141259 290175
rect 140949 290113 141259 290147
rect 140949 290085 140997 290113
rect 141025 290085 141059 290113
rect 141087 290085 141121 290113
rect 141149 290085 141183 290113
rect 141211 290085 141259 290113
rect 140949 290051 141259 290085
rect 140949 290023 140997 290051
rect 141025 290023 141059 290051
rect 141087 290023 141121 290051
rect 141149 290023 141183 290051
rect 141211 290023 141259 290051
rect 140949 289989 141259 290023
rect 140949 289961 140997 289989
rect 141025 289961 141059 289989
rect 141087 289961 141121 289989
rect 141149 289961 141183 289989
rect 141211 289961 141259 289989
rect 140949 281175 141259 289961
rect 140949 281147 140997 281175
rect 141025 281147 141059 281175
rect 141087 281147 141121 281175
rect 141149 281147 141183 281175
rect 141211 281147 141259 281175
rect 140949 281113 141259 281147
rect 140949 281085 140997 281113
rect 141025 281085 141059 281113
rect 141087 281085 141121 281113
rect 141149 281085 141183 281113
rect 141211 281085 141259 281113
rect 140949 281051 141259 281085
rect 140949 281023 140997 281051
rect 141025 281023 141059 281051
rect 141087 281023 141121 281051
rect 141149 281023 141183 281051
rect 141211 281023 141259 281051
rect 140949 280989 141259 281023
rect 140949 280961 140997 280989
rect 141025 280961 141059 280989
rect 141087 280961 141121 280989
rect 141149 280961 141183 280989
rect 141211 280961 141259 280989
rect 140949 272175 141259 280961
rect 140949 272147 140997 272175
rect 141025 272147 141059 272175
rect 141087 272147 141121 272175
rect 141149 272147 141183 272175
rect 141211 272147 141259 272175
rect 140949 272113 141259 272147
rect 140949 272085 140997 272113
rect 141025 272085 141059 272113
rect 141087 272085 141121 272113
rect 141149 272085 141183 272113
rect 141211 272085 141259 272113
rect 140949 272051 141259 272085
rect 140949 272023 140997 272051
rect 141025 272023 141059 272051
rect 141087 272023 141121 272051
rect 141149 272023 141183 272051
rect 141211 272023 141259 272051
rect 140949 271989 141259 272023
rect 140949 271961 140997 271989
rect 141025 271961 141059 271989
rect 141087 271961 141121 271989
rect 141149 271961 141183 271989
rect 141211 271961 141259 271989
rect 140949 268935 141259 271961
rect 142809 299086 143119 299134
rect 142809 299058 142857 299086
rect 142885 299058 142919 299086
rect 142947 299058 142981 299086
rect 143009 299058 143043 299086
rect 143071 299058 143119 299086
rect 142809 299024 143119 299058
rect 142809 298996 142857 299024
rect 142885 298996 142919 299024
rect 142947 298996 142981 299024
rect 143009 298996 143043 299024
rect 143071 298996 143119 299024
rect 142809 298962 143119 298996
rect 142809 298934 142857 298962
rect 142885 298934 142919 298962
rect 142947 298934 142981 298962
rect 143009 298934 143043 298962
rect 143071 298934 143119 298962
rect 142809 298900 143119 298934
rect 142809 298872 142857 298900
rect 142885 298872 142919 298900
rect 142947 298872 142981 298900
rect 143009 298872 143043 298900
rect 143071 298872 143119 298900
rect 142809 293175 143119 298872
rect 142809 293147 142857 293175
rect 142885 293147 142919 293175
rect 142947 293147 142981 293175
rect 143009 293147 143043 293175
rect 143071 293147 143119 293175
rect 142809 293113 143119 293147
rect 142809 293085 142857 293113
rect 142885 293085 142919 293113
rect 142947 293085 142981 293113
rect 143009 293085 143043 293113
rect 143071 293085 143119 293113
rect 142809 293051 143119 293085
rect 142809 293023 142857 293051
rect 142885 293023 142919 293051
rect 142947 293023 142981 293051
rect 143009 293023 143043 293051
rect 143071 293023 143119 293051
rect 142809 292989 143119 293023
rect 142809 292961 142857 292989
rect 142885 292961 142919 292989
rect 142947 292961 142981 292989
rect 143009 292961 143043 292989
rect 143071 292961 143119 292989
rect 142809 284175 143119 292961
rect 142809 284147 142857 284175
rect 142885 284147 142919 284175
rect 142947 284147 142981 284175
rect 143009 284147 143043 284175
rect 143071 284147 143119 284175
rect 142809 284113 143119 284147
rect 142809 284085 142857 284113
rect 142885 284085 142919 284113
rect 142947 284085 142981 284113
rect 143009 284085 143043 284113
rect 143071 284085 143119 284113
rect 142809 284051 143119 284085
rect 142809 284023 142857 284051
rect 142885 284023 142919 284051
rect 142947 284023 142981 284051
rect 143009 284023 143043 284051
rect 143071 284023 143119 284051
rect 142809 283989 143119 284023
rect 142809 283961 142857 283989
rect 142885 283961 142919 283989
rect 142947 283961 142981 283989
rect 143009 283961 143043 283989
rect 143071 283961 143119 283989
rect 142809 275175 143119 283961
rect 142809 275147 142857 275175
rect 142885 275147 142919 275175
rect 142947 275147 142981 275175
rect 143009 275147 143043 275175
rect 143071 275147 143119 275175
rect 142809 275113 143119 275147
rect 142809 275085 142857 275113
rect 142885 275085 142919 275113
rect 142947 275085 142981 275113
rect 143009 275085 143043 275113
rect 143071 275085 143119 275113
rect 142809 275051 143119 275085
rect 142809 275023 142857 275051
rect 142885 275023 142919 275051
rect 142947 275023 142981 275051
rect 143009 275023 143043 275051
rect 143071 275023 143119 275051
rect 142809 274989 143119 275023
rect 142809 274961 142857 274989
rect 142885 274961 142919 274989
rect 142947 274961 142981 274989
rect 143009 274961 143043 274989
rect 143071 274961 143119 274989
rect 142809 268935 143119 274961
rect 156309 298606 156619 299134
rect 156309 298578 156357 298606
rect 156385 298578 156419 298606
rect 156447 298578 156481 298606
rect 156509 298578 156543 298606
rect 156571 298578 156619 298606
rect 156309 298544 156619 298578
rect 156309 298516 156357 298544
rect 156385 298516 156419 298544
rect 156447 298516 156481 298544
rect 156509 298516 156543 298544
rect 156571 298516 156619 298544
rect 156309 298482 156619 298516
rect 156309 298454 156357 298482
rect 156385 298454 156419 298482
rect 156447 298454 156481 298482
rect 156509 298454 156543 298482
rect 156571 298454 156619 298482
rect 156309 298420 156619 298454
rect 156309 298392 156357 298420
rect 156385 298392 156419 298420
rect 156447 298392 156481 298420
rect 156509 298392 156543 298420
rect 156571 298392 156619 298420
rect 156309 290175 156619 298392
rect 156309 290147 156357 290175
rect 156385 290147 156419 290175
rect 156447 290147 156481 290175
rect 156509 290147 156543 290175
rect 156571 290147 156619 290175
rect 156309 290113 156619 290147
rect 156309 290085 156357 290113
rect 156385 290085 156419 290113
rect 156447 290085 156481 290113
rect 156509 290085 156543 290113
rect 156571 290085 156619 290113
rect 156309 290051 156619 290085
rect 156309 290023 156357 290051
rect 156385 290023 156419 290051
rect 156447 290023 156481 290051
rect 156509 290023 156543 290051
rect 156571 290023 156619 290051
rect 156309 289989 156619 290023
rect 156309 289961 156357 289989
rect 156385 289961 156419 289989
rect 156447 289961 156481 289989
rect 156509 289961 156543 289989
rect 156571 289961 156619 289989
rect 156309 281175 156619 289961
rect 156309 281147 156357 281175
rect 156385 281147 156419 281175
rect 156447 281147 156481 281175
rect 156509 281147 156543 281175
rect 156571 281147 156619 281175
rect 156309 281113 156619 281147
rect 156309 281085 156357 281113
rect 156385 281085 156419 281113
rect 156447 281085 156481 281113
rect 156509 281085 156543 281113
rect 156571 281085 156619 281113
rect 156309 281051 156619 281085
rect 156309 281023 156357 281051
rect 156385 281023 156419 281051
rect 156447 281023 156481 281051
rect 156509 281023 156543 281051
rect 156571 281023 156619 281051
rect 156309 280989 156619 281023
rect 156309 280961 156357 280989
rect 156385 280961 156419 280989
rect 156447 280961 156481 280989
rect 156509 280961 156543 280989
rect 156571 280961 156619 280989
rect 156309 272175 156619 280961
rect 156309 272147 156357 272175
rect 156385 272147 156419 272175
rect 156447 272147 156481 272175
rect 156509 272147 156543 272175
rect 156571 272147 156619 272175
rect 156309 272113 156619 272147
rect 156309 272085 156357 272113
rect 156385 272085 156419 272113
rect 156447 272085 156481 272113
rect 156509 272085 156543 272113
rect 156571 272085 156619 272113
rect 156309 272051 156619 272085
rect 156309 272023 156357 272051
rect 156385 272023 156419 272051
rect 156447 272023 156481 272051
rect 156509 272023 156543 272051
rect 156571 272023 156619 272051
rect 156309 271989 156619 272023
rect 156309 271961 156357 271989
rect 156385 271961 156419 271989
rect 156447 271961 156481 271989
rect 156509 271961 156543 271989
rect 156571 271961 156619 271989
rect 156309 268935 156619 271961
rect 158169 299086 158479 299134
rect 158169 299058 158217 299086
rect 158245 299058 158279 299086
rect 158307 299058 158341 299086
rect 158369 299058 158403 299086
rect 158431 299058 158479 299086
rect 158169 299024 158479 299058
rect 158169 298996 158217 299024
rect 158245 298996 158279 299024
rect 158307 298996 158341 299024
rect 158369 298996 158403 299024
rect 158431 298996 158479 299024
rect 158169 298962 158479 298996
rect 158169 298934 158217 298962
rect 158245 298934 158279 298962
rect 158307 298934 158341 298962
rect 158369 298934 158403 298962
rect 158431 298934 158479 298962
rect 158169 298900 158479 298934
rect 158169 298872 158217 298900
rect 158245 298872 158279 298900
rect 158307 298872 158341 298900
rect 158369 298872 158403 298900
rect 158431 298872 158479 298900
rect 158169 293175 158479 298872
rect 158169 293147 158217 293175
rect 158245 293147 158279 293175
rect 158307 293147 158341 293175
rect 158369 293147 158403 293175
rect 158431 293147 158479 293175
rect 158169 293113 158479 293147
rect 158169 293085 158217 293113
rect 158245 293085 158279 293113
rect 158307 293085 158341 293113
rect 158369 293085 158403 293113
rect 158431 293085 158479 293113
rect 158169 293051 158479 293085
rect 158169 293023 158217 293051
rect 158245 293023 158279 293051
rect 158307 293023 158341 293051
rect 158369 293023 158403 293051
rect 158431 293023 158479 293051
rect 158169 292989 158479 293023
rect 158169 292961 158217 292989
rect 158245 292961 158279 292989
rect 158307 292961 158341 292989
rect 158369 292961 158403 292989
rect 158431 292961 158479 292989
rect 158169 284175 158479 292961
rect 158169 284147 158217 284175
rect 158245 284147 158279 284175
rect 158307 284147 158341 284175
rect 158369 284147 158403 284175
rect 158431 284147 158479 284175
rect 158169 284113 158479 284147
rect 158169 284085 158217 284113
rect 158245 284085 158279 284113
rect 158307 284085 158341 284113
rect 158369 284085 158403 284113
rect 158431 284085 158479 284113
rect 158169 284051 158479 284085
rect 158169 284023 158217 284051
rect 158245 284023 158279 284051
rect 158307 284023 158341 284051
rect 158369 284023 158403 284051
rect 158431 284023 158479 284051
rect 158169 283989 158479 284023
rect 158169 283961 158217 283989
rect 158245 283961 158279 283989
rect 158307 283961 158341 283989
rect 158369 283961 158403 283989
rect 158431 283961 158479 283989
rect 158169 275175 158479 283961
rect 158169 275147 158217 275175
rect 158245 275147 158279 275175
rect 158307 275147 158341 275175
rect 158369 275147 158403 275175
rect 158431 275147 158479 275175
rect 158169 275113 158479 275147
rect 158169 275085 158217 275113
rect 158245 275085 158279 275113
rect 158307 275085 158341 275113
rect 158369 275085 158403 275113
rect 158431 275085 158479 275113
rect 158169 275051 158479 275085
rect 158169 275023 158217 275051
rect 158245 275023 158279 275051
rect 158307 275023 158341 275051
rect 158369 275023 158403 275051
rect 158431 275023 158479 275051
rect 158169 274989 158479 275023
rect 158169 274961 158217 274989
rect 158245 274961 158279 274989
rect 158307 274961 158341 274989
rect 158369 274961 158403 274989
rect 158431 274961 158479 274989
rect 158169 268935 158479 274961
rect 171669 298606 171979 299134
rect 171669 298578 171717 298606
rect 171745 298578 171779 298606
rect 171807 298578 171841 298606
rect 171869 298578 171903 298606
rect 171931 298578 171979 298606
rect 171669 298544 171979 298578
rect 171669 298516 171717 298544
rect 171745 298516 171779 298544
rect 171807 298516 171841 298544
rect 171869 298516 171903 298544
rect 171931 298516 171979 298544
rect 171669 298482 171979 298516
rect 171669 298454 171717 298482
rect 171745 298454 171779 298482
rect 171807 298454 171841 298482
rect 171869 298454 171903 298482
rect 171931 298454 171979 298482
rect 171669 298420 171979 298454
rect 171669 298392 171717 298420
rect 171745 298392 171779 298420
rect 171807 298392 171841 298420
rect 171869 298392 171903 298420
rect 171931 298392 171979 298420
rect 171669 290175 171979 298392
rect 171669 290147 171717 290175
rect 171745 290147 171779 290175
rect 171807 290147 171841 290175
rect 171869 290147 171903 290175
rect 171931 290147 171979 290175
rect 171669 290113 171979 290147
rect 171669 290085 171717 290113
rect 171745 290085 171779 290113
rect 171807 290085 171841 290113
rect 171869 290085 171903 290113
rect 171931 290085 171979 290113
rect 171669 290051 171979 290085
rect 171669 290023 171717 290051
rect 171745 290023 171779 290051
rect 171807 290023 171841 290051
rect 171869 290023 171903 290051
rect 171931 290023 171979 290051
rect 171669 289989 171979 290023
rect 171669 289961 171717 289989
rect 171745 289961 171779 289989
rect 171807 289961 171841 289989
rect 171869 289961 171903 289989
rect 171931 289961 171979 289989
rect 171669 281175 171979 289961
rect 171669 281147 171717 281175
rect 171745 281147 171779 281175
rect 171807 281147 171841 281175
rect 171869 281147 171903 281175
rect 171931 281147 171979 281175
rect 171669 281113 171979 281147
rect 171669 281085 171717 281113
rect 171745 281085 171779 281113
rect 171807 281085 171841 281113
rect 171869 281085 171903 281113
rect 171931 281085 171979 281113
rect 171669 281051 171979 281085
rect 171669 281023 171717 281051
rect 171745 281023 171779 281051
rect 171807 281023 171841 281051
rect 171869 281023 171903 281051
rect 171931 281023 171979 281051
rect 171669 280989 171979 281023
rect 171669 280961 171717 280989
rect 171745 280961 171779 280989
rect 171807 280961 171841 280989
rect 171869 280961 171903 280989
rect 171931 280961 171979 280989
rect 171669 272175 171979 280961
rect 171669 272147 171717 272175
rect 171745 272147 171779 272175
rect 171807 272147 171841 272175
rect 171869 272147 171903 272175
rect 171931 272147 171979 272175
rect 171669 272113 171979 272147
rect 171669 272085 171717 272113
rect 171745 272085 171779 272113
rect 171807 272085 171841 272113
rect 171869 272085 171903 272113
rect 171931 272085 171979 272113
rect 171669 272051 171979 272085
rect 171669 272023 171717 272051
rect 171745 272023 171779 272051
rect 171807 272023 171841 272051
rect 171869 272023 171903 272051
rect 171931 272023 171979 272051
rect 171669 271989 171979 272023
rect 171669 271961 171717 271989
rect 171745 271961 171779 271989
rect 171807 271961 171841 271989
rect 171869 271961 171903 271989
rect 171931 271961 171979 271989
rect 96729 266147 96777 266175
rect 96805 266147 96839 266175
rect 96867 266147 96901 266175
rect 96929 266147 96963 266175
rect 96991 266147 97039 266175
rect 96729 266113 97039 266147
rect 96729 266085 96777 266113
rect 96805 266085 96839 266113
rect 96867 266085 96901 266113
rect 96929 266085 96963 266113
rect 96991 266085 97039 266113
rect 96729 266051 97039 266085
rect 96729 266023 96777 266051
rect 96805 266023 96839 266051
rect 96867 266023 96901 266051
rect 96929 266023 96963 266051
rect 96991 266023 97039 266051
rect 96729 265989 97039 266023
rect 96729 265961 96777 265989
rect 96805 265961 96839 265989
rect 96867 265961 96901 265989
rect 96929 265961 96963 265989
rect 96991 265961 97039 265989
rect 96729 257175 97039 265961
rect 109904 266175 110064 266192
rect 109904 266147 109939 266175
rect 109967 266147 110001 266175
rect 110029 266147 110064 266175
rect 109904 266113 110064 266147
rect 109904 266085 109939 266113
rect 109967 266085 110001 266113
rect 110029 266085 110064 266113
rect 109904 266051 110064 266085
rect 109904 266023 109939 266051
rect 109967 266023 110001 266051
rect 110029 266023 110064 266051
rect 109904 265989 110064 266023
rect 109904 265961 109939 265989
rect 109967 265961 110001 265989
rect 110029 265961 110064 265989
rect 109904 265944 110064 265961
rect 125264 266175 125424 266192
rect 125264 266147 125299 266175
rect 125327 266147 125361 266175
rect 125389 266147 125424 266175
rect 125264 266113 125424 266147
rect 125264 266085 125299 266113
rect 125327 266085 125361 266113
rect 125389 266085 125424 266113
rect 125264 266051 125424 266085
rect 125264 266023 125299 266051
rect 125327 266023 125361 266051
rect 125389 266023 125424 266051
rect 125264 265989 125424 266023
rect 125264 265961 125299 265989
rect 125327 265961 125361 265989
rect 125389 265961 125424 265989
rect 125264 265944 125424 265961
rect 140624 266175 140784 266192
rect 140624 266147 140659 266175
rect 140687 266147 140721 266175
rect 140749 266147 140784 266175
rect 140624 266113 140784 266147
rect 140624 266085 140659 266113
rect 140687 266085 140721 266113
rect 140749 266085 140784 266113
rect 140624 266051 140784 266085
rect 140624 266023 140659 266051
rect 140687 266023 140721 266051
rect 140749 266023 140784 266051
rect 140624 265989 140784 266023
rect 140624 265961 140659 265989
rect 140687 265961 140721 265989
rect 140749 265961 140784 265989
rect 140624 265944 140784 265961
rect 155984 266175 156144 266192
rect 155984 266147 156019 266175
rect 156047 266147 156081 266175
rect 156109 266147 156144 266175
rect 155984 266113 156144 266147
rect 155984 266085 156019 266113
rect 156047 266085 156081 266113
rect 156109 266085 156144 266113
rect 155984 266051 156144 266085
rect 155984 266023 156019 266051
rect 156047 266023 156081 266051
rect 156109 266023 156144 266051
rect 155984 265989 156144 266023
rect 155984 265961 156019 265989
rect 156047 265961 156081 265989
rect 156109 265961 156144 265989
rect 155984 265944 156144 265961
rect 102224 263175 102384 263192
rect 102224 263147 102259 263175
rect 102287 263147 102321 263175
rect 102349 263147 102384 263175
rect 102224 263113 102384 263147
rect 102224 263085 102259 263113
rect 102287 263085 102321 263113
rect 102349 263085 102384 263113
rect 102224 263051 102384 263085
rect 102224 263023 102259 263051
rect 102287 263023 102321 263051
rect 102349 263023 102384 263051
rect 102224 262989 102384 263023
rect 102224 262961 102259 262989
rect 102287 262961 102321 262989
rect 102349 262961 102384 262989
rect 102224 262944 102384 262961
rect 117584 263175 117744 263192
rect 117584 263147 117619 263175
rect 117647 263147 117681 263175
rect 117709 263147 117744 263175
rect 117584 263113 117744 263147
rect 117584 263085 117619 263113
rect 117647 263085 117681 263113
rect 117709 263085 117744 263113
rect 117584 263051 117744 263085
rect 117584 263023 117619 263051
rect 117647 263023 117681 263051
rect 117709 263023 117744 263051
rect 117584 262989 117744 263023
rect 117584 262961 117619 262989
rect 117647 262961 117681 262989
rect 117709 262961 117744 262989
rect 117584 262944 117744 262961
rect 132944 263175 133104 263192
rect 132944 263147 132979 263175
rect 133007 263147 133041 263175
rect 133069 263147 133104 263175
rect 132944 263113 133104 263147
rect 132944 263085 132979 263113
rect 133007 263085 133041 263113
rect 133069 263085 133104 263113
rect 132944 263051 133104 263085
rect 132944 263023 132979 263051
rect 133007 263023 133041 263051
rect 133069 263023 133104 263051
rect 132944 262989 133104 263023
rect 132944 262961 132979 262989
rect 133007 262961 133041 262989
rect 133069 262961 133104 262989
rect 132944 262944 133104 262961
rect 148304 263175 148464 263192
rect 148304 263147 148339 263175
rect 148367 263147 148401 263175
rect 148429 263147 148464 263175
rect 148304 263113 148464 263147
rect 148304 263085 148339 263113
rect 148367 263085 148401 263113
rect 148429 263085 148464 263113
rect 148304 263051 148464 263085
rect 148304 263023 148339 263051
rect 148367 263023 148401 263051
rect 148429 263023 148464 263051
rect 148304 262989 148464 263023
rect 148304 262961 148339 262989
rect 148367 262961 148401 262989
rect 148429 262961 148464 262989
rect 148304 262944 148464 262961
rect 163664 263175 163824 263192
rect 163664 263147 163699 263175
rect 163727 263147 163761 263175
rect 163789 263147 163824 263175
rect 163664 263113 163824 263147
rect 163664 263085 163699 263113
rect 163727 263085 163761 263113
rect 163789 263085 163824 263113
rect 163664 263051 163824 263085
rect 163664 263023 163699 263051
rect 163727 263023 163761 263051
rect 163789 263023 163824 263051
rect 163664 262989 163824 263023
rect 163664 262961 163699 262989
rect 163727 262961 163761 262989
rect 163789 262961 163824 262989
rect 163664 262944 163824 262961
rect 171669 263175 171979 271961
rect 171669 263147 171717 263175
rect 171745 263147 171779 263175
rect 171807 263147 171841 263175
rect 171869 263147 171903 263175
rect 171931 263147 171979 263175
rect 171669 263113 171979 263147
rect 171669 263085 171717 263113
rect 171745 263085 171779 263113
rect 171807 263085 171841 263113
rect 171869 263085 171903 263113
rect 171931 263085 171979 263113
rect 171669 263051 171979 263085
rect 171669 263023 171717 263051
rect 171745 263023 171779 263051
rect 171807 263023 171841 263051
rect 171869 263023 171903 263051
rect 171931 263023 171979 263051
rect 171669 262989 171979 263023
rect 171669 262961 171717 262989
rect 171745 262961 171779 262989
rect 171807 262961 171841 262989
rect 171869 262961 171903 262989
rect 171931 262961 171979 262989
rect 96729 257147 96777 257175
rect 96805 257147 96839 257175
rect 96867 257147 96901 257175
rect 96929 257147 96963 257175
rect 96991 257147 97039 257175
rect 96729 257113 97039 257147
rect 96729 257085 96777 257113
rect 96805 257085 96839 257113
rect 96867 257085 96901 257113
rect 96929 257085 96963 257113
rect 96991 257085 97039 257113
rect 96729 257051 97039 257085
rect 96729 257023 96777 257051
rect 96805 257023 96839 257051
rect 96867 257023 96901 257051
rect 96929 257023 96963 257051
rect 96991 257023 97039 257051
rect 96729 256989 97039 257023
rect 96729 256961 96777 256989
rect 96805 256961 96839 256989
rect 96867 256961 96901 256989
rect 96929 256961 96963 256989
rect 96991 256961 97039 256989
rect 96729 248175 97039 256961
rect 109904 257175 110064 257192
rect 109904 257147 109939 257175
rect 109967 257147 110001 257175
rect 110029 257147 110064 257175
rect 109904 257113 110064 257147
rect 109904 257085 109939 257113
rect 109967 257085 110001 257113
rect 110029 257085 110064 257113
rect 109904 257051 110064 257085
rect 109904 257023 109939 257051
rect 109967 257023 110001 257051
rect 110029 257023 110064 257051
rect 109904 256989 110064 257023
rect 109904 256961 109939 256989
rect 109967 256961 110001 256989
rect 110029 256961 110064 256989
rect 109904 256944 110064 256961
rect 125264 257175 125424 257192
rect 125264 257147 125299 257175
rect 125327 257147 125361 257175
rect 125389 257147 125424 257175
rect 125264 257113 125424 257147
rect 125264 257085 125299 257113
rect 125327 257085 125361 257113
rect 125389 257085 125424 257113
rect 125264 257051 125424 257085
rect 125264 257023 125299 257051
rect 125327 257023 125361 257051
rect 125389 257023 125424 257051
rect 125264 256989 125424 257023
rect 125264 256961 125299 256989
rect 125327 256961 125361 256989
rect 125389 256961 125424 256989
rect 125264 256944 125424 256961
rect 140624 257175 140784 257192
rect 140624 257147 140659 257175
rect 140687 257147 140721 257175
rect 140749 257147 140784 257175
rect 140624 257113 140784 257147
rect 140624 257085 140659 257113
rect 140687 257085 140721 257113
rect 140749 257085 140784 257113
rect 140624 257051 140784 257085
rect 140624 257023 140659 257051
rect 140687 257023 140721 257051
rect 140749 257023 140784 257051
rect 140624 256989 140784 257023
rect 140624 256961 140659 256989
rect 140687 256961 140721 256989
rect 140749 256961 140784 256989
rect 140624 256944 140784 256961
rect 155984 257175 156144 257192
rect 155984 257147 156019 257175
rect 156047 257147 156081 257175
rect 156109 257147 156144 257175
rect 155984 257113 156144 257147
rect 155984 257085 156019 257113
rect 156047 257085 156081 257113
rect 156109 257085 156144 257113
rect 155984 257051 156144 257085
rect 155984 257023 156019 257051
rect 156047 257023 156081 257051
rect 156109 257023 156144 257051
rect 155984 256989 156144 257023
rect 155984 256961 156019 256989
rect 156047 256961 156081 256989
rect 156109 256961 156144 256989
rect 155984 256944 156144 256961
rect 102224 254175 102384 254192
rect 102224 254147 102259 254175
rect 102287 254147 102321 254175
rect 102349 254147 102384 254175
rect 102224 254113 102384 254147
rect 102224 254085 102259 254113
rect 102287 254085 102321 254113
rect 102349 254085 102384 254113
rect 102224 254051 102384 254085
rect 102224 254023 102259 254051
rect 102287 254023 102321 254051
rect 102349 254023 102384 254051
rect 102224 253989 102384 254023
rect 102224 253961 102259 253989
rect 102287 253961 102321 253989
rect 102349 253961 102384 253989
rect 102224 253944 102384 253961
rect 117584 254175 117744 254192
rect 117584 254147 117619 254175
rect 117647 254147 117681 254175
rect 117709 254147 117744 254175
rect 117584 254113 117744 254147
rect 117584 254085 117619 254113
rect 117647 254085 117681 254113
rect 117709 254085 117744 254113
rect 117584 254051 117744 254085
rect 117584 254023 117619 254051
rect 117647 254023 117681 254051
rect 117709 254023 117744 254051
rect 117584 253989 117744 254023
rect 117584 253961 117619 253989
rect 117647 253961 117681 253989
rect 117709 253961 117744 253989
rect 117584 253944 117744 253961
rect 132944 254175 133104 254192
rect 132944 254147 132979 254175
rect 133007 254147 133041 254175
rect 133069 254147 133104 254175
rect 132944 254113 133104 254147
rect 132944 254085 132979 254113
rect 133007 254085 133041 254113
rect 133069 254085 133104 254113
rect 132944 254051 133104 254085
rect 132944 254023 132979 254051
rect 133007 254023 133041 254051
rect 133069 254023 133104 254051
rect 132944 253989 133104 254023
rect 132944 253961 132979 253989
rect 133007 253961 133041 253989
rect 133069 253961 133104 253989
rect 132944 253944 133104 253961
rect 148304 254175 148464 254192
rect 148304 254147 148339 254175
rect 148367 254147 148401 254175
rect 148429 254147 148464 254175
rect 148304 254113 148464 254147
rect 148304 254085 148339 254113
rect 148367 254085 148401 254113
rect 148429 254085 148464 254113
rect 148304 254051 148464 254085
rect 148304 254023 148339 254051
rect 148367 254023 148401 254051
rect 148429 254023 148464 254051
rect 148304 253989 148464 254023
rect 148304 253961 148339 253989
rect 148367 253961 148401 253989
rect 148429 253961 148464 253989
rect 148304 253944 148464 253961
rect 163664 254175 163824 254192
rect 163664 254147 163699 254175
rect 163727 254147 163761 254175
rect 163789 254147 163824 254175
rect 163664 254113 163824 254147
rect 163664 254085 163699 254113
rect 163727 254085 163761 254113
rect 163789 254085 163824 254113
rect 163664 254051 163824 254085
rect 163664 254023 163699 254051
rect 163727 254023 163761 254051
rect 163789 254023 163824 254051
rect 163664 253989 163824 254023
rect 163664 253961 163699 253989
rect 163727 253961 163761 253989
rect 163789 253961 163824 253989
rect 163664 253944 163824 253961
rect 171669 254175 171979 262961
rect 171669 254147 171717 254175
rect 171745 254147 171779 254175
rect 171807 254147 171841 254175
rect 171869 254147 171903 254175
rect 171931 254147 171979 254175
rect 171669 254113 171979 254147
rect 171669 254085 171717 254113
rect 171745 254085 171779 254113
rect 171807 254085 171841 254113
rect 171869 254085 171903 254113
rect 171931 254085 171979 254113
rect 171669 254051 171979 254085
rect 171669 254023 171717 254051
rect 171745 254023 171779 254051
rect 171807 254023 171841 254051
rect 171869 254023 171903 254051
rect 171931 254023 171979 254051
rect 171669 253989 171979 254023
rect 171669 253961 171717 253989
rect 171745 253961 171779 253989
rect 171807 253961 171841 253989
rect 171869 253961 171903 253989
rect 171931 253961 171979 253989
rect 96729 248147 96777 248175
rect 96805 248147 96839 248175
rect 96867 248147 96901 248175
rect 96929 248147 96963 248175
rect 96991 248147 97039 248175
rect 96729 248113 97039 248147
rect 96729 248085 96777 248113
rect 96805 248085 96839 248113
rect 96867 248085 96901 248113
rect 96929 248085 96963 248113
rect 96991 248085 97039 248113
rect 96729 248051 97039 248085
rect 96729 248023 96777 248051
rect 96805 248023 96839 248051
rect 96867 248023 96901 248051
rect 96929 248023 96963 248051
rect 96991 248023 97039 248051
rect 96729 247989 97039 248023
rect 96729 247961 96777 247989
rect 96805 247961 96839 247989
rect 96867 247961 96901 247989
rect 96929 247961 96963 247989
rect 96991 247961 97039 247989
rect 96729 239175 97039 247961
rect 109904 248175 110064 248192
rect 109904 248147 109939 248175
rect 109967 248147 110001 248175
rect 110029 248147 110064 248175
rect 109904 248113 110064 248147
rect 109904 248085 109939 248113
rect 109967 248085 110001 248113
rect 110029 248085 110064 248113
rect 109904 248051 110064 248085
rect 109904 248023 109939 248051
rect 109967 248023 110001 248051
rect 110029 248023 110064 248051
rect 109904 247989 110064 248023
rect 109904 247961 109939 247989
rect 109967 247961 110001 247989
rect 110029 247961 110064 247989
rect 109904 247944 110064 247961
rect 125264 248175 125424 248192
rect 125264 248147 125299 248175
rect 125327 248147 125361 248175
rect 125389 248147 125424 248175
rect 125264 248113 125424 248147
rect 125264 248085 125299 248113
rect 125327 248085 125361 248113
rect 125389 248085 125424 248113
rect 125264 248051 125424 248085
rect 125264 248023 125299 248051
rect 125327 248023 125361 248051
rect 125389 248023 125424 248051
rect 125264 247989 125424 248023
rect 125264 247961 125299 247989
rect 125327 247961 125361 247989
rect 125389 247961 125424 247989
rect 125264 247944 125424 247961
rect 140624 248175 140784 248192
rect 140624 248147 140659 248175
rect 140687 248147 140721 248175
rect 140749 248147 140784 248175
rect 140624 248113 140784 248147
rect 140624 248085 140659 248113
rect 140687 248085 140721 248113
rect 140749 248085 140784 248113
rect 140624 248051 140784 248085
rect 140624 248023 140659 248051
rect 140687 248023 140721 248051
rect 140749 248023 140784 248051
rect 140624 247989 140784 248023
rect 140624 247961 140659 247989
rect 140687 247961 140721 247989
rect 140749 247961 140784 247989
rect 140624 247944 140784 247961
rect 155984 248175 156144 248192
rect 155984 248147 156019 248175
rect 156047 248147 156081 248175
rect 156109 248147 156144 248175
rect 155984 248113 156144 248147
rect 155984 248085 156019 248113
rect 156047 248085 156081 248113
rect 156109 248085 156144 248113
rect 155984 248051 156144 248085
rect 155984 248023 156019 248051
rect 156047 248023 156081 248051
rect 156109 248023 156144 248051
rect 155984 247989 156144 248023
rect 155984 247961 156019 247989
rect 156047 247961 156081 247989
rect 156109 247961 156144 247989
rect 155984 247944 156144 247961
rect 102224 245175 102384 245192
rect 102224 245147 102259 245175
rect 102287 245147 102321 245175
rect 102349 245147 102384 245175
rect 102224 245113 102384 245147
rect 102224 245085 102259 245113
rect 102287 245085 102321 245113
rect 102349 245085 102384 245113
rect 102224 245051 102384 245085
rect 102224 245023 102259 245051
rect 102287 245023 102321 245051
rect 102349 245023 102384 245051
rect 102224 244989 102384 245023
rect 102224 244961 102259 244989
rect 102287 244961 102321 244989
rect 102349 244961 102384 244989
rect 102224 244944 102384 244961
rect 117584 245175 117744 245192
rect 117584 245147 117619 245175
rect 117647 245147 117681 245175
rect 117709 245147 117744 245175
rect 117584 245113 117744 245147
rect 117584 245085 117619 245113
rect 117647 245085 117681 245113
rect 117709 245085 117744 245113
rect 117584 245051 117744 245085
rect 117584 245023 117619 245051
rect 117647 245023 117681 245051
rect 117709 245023 117744 245051
rect 117584 244989 117744 245023
rect 117584 244961 117619 244989
rect 117647 244961 117681 244989
rect 117709 244961 117744 244989
rect 117584 244944 117744 244961
rect 132944 245175 133104 245192
rect 132944 245147 132979 245175
rect 133007 245147 133041 245175
rect 133069 245147 133104 245175
rect 132944 245113 133104 245147
rect 132944 245085 132979 245113
rect 133007 245085 133041 245113
rect 133069 245085 133104 245113
rect 132944 245051 133104 245085
rect 132944 245023 132979 245051
rect 133007 245023 133041 245051
rect 133069 245023 133104 245051
rect 132944 244989 133104 245023
rect 132944 244961 132979 244989
rect 133007 244961 133041 244989
rect 133069 244961 133104 244989
rect 132944 244944 133104 244961
rect 148304 245175 148464 245192
rect 148304 245147 148339 245175
rect 148367 245147 148401 245175
rect 148429 245147 148464 245175
rect 148304 245113 148464 245147
rect 148304 245085 148339 245113
rect 148367 245085 148401 245113
rect 148429 245085 148464 245113
rect 148304 245051 148464 245085
rect 148304 245023 148339 245051
rect 148367 245023 148401 245051
rect 148429 245023 148464 245051
rect 148304 244989 148464 245023
rect 148304 244961 148339 244989
rect 148367 244961 148401 244989
rect 148429 244961 148464 244989
rect 148304 244944 148464 244961
rect 163664 245175 163824 245192
rect 163664 245147 163699 245175
rect 163727 245147 163761 245175
rect 163789 245147 163824 245175
rect 163664 245113 163824 245147
rect 163664 245085 163699 245113
rect 163727 245085 163761 245113
rect 163789 245085 163824 245113
rect 163664 245051 163824 245085
rect 163664 245023 163699 245051
rect 163727 245023 163761 245051
rect 163789 245023 163824 245051
rect 163664 244989 163824 245023
rect 163664 244961 163699 244989
rect 163727 244961 163761 244989
rect 163789 244961 163824 244989
rect 163664 244944 163824 244961
rect 171669 245175 171979 253961
rect 171669 245147 171717 245175
rect 171745 245147 171779 245175
rect 171807 245147 171841 245175
rect 171869 245147 171903 245175
rect 171931 245147 171979 245175
rect 171669 245113 171979 245147
rect 171669 245085 171717 245113
rect 171745 245085 171779 245113
rect 171807 245085 171841 245113
rect 171869 245085 171903 245113
rect 171931 245085 171979 245113
rect 171669 245051 171979 245085
rect 171669 245023 171717 245051
rect 171745 245023 171779 245051
rect 171807 245023 171841 245051
rect 171869 245023 171903 245051
rect 171931 245023 171979 245051
rect 171669 244989 171979 245023
rect 171669 244961 171717 244989
rect 171745 244961 171779 244989
rect 171807 244961 171841 244989
rect 171869 244961 171903 244989
rect 171931 244961 171979 244989
rect 96729 239147 96777 239175
rect 96805 239147 96839 239175
rect 96867 239147 96901 239175
rect 96929 239147 96963 239175
rect 96991 239147 97039 239175
rect 96729 239113 97039 239147
rect 96729 239085 96777 239113
rect 96805 239085 96839 239113
rect 96867 239085 96901 239113
rect 96929 239085 96963 239113
rect 96991 239085 97039 239113
rect 96729 239051 97039 239085
rect 96729 239023 96777 239051
rect 96805 239023 96839 239051
rect 96867 239023 96901 239051
rect 96929 239023 96963 239051
rect 96991 239023 97039 239051
rect 96729 238989 97039 239023
rect 96729 238961 96777 238989
rect 96805 238961 96839 238989
rect 96867 238961 96901 238989
rect 96929 238961 96963 238989
rect 96991 238961 97039 238989
rect 96729 230175 97039 238961
rect 109904 239175 110064 239192
rect 109904 239147 109939 239175
rect 109967 239147 110001 239175
rect 110029 239147 110064 239175
rect 109904 239113 110064 239147
rect 109904 239085 109939 239113
rect 109967 239085 110001 239113
rect 110029 239085 110064 239113
rect 109904 239051 110064 239085
rect 109904 239023 109939 239051
rect 109967 239023 110001 239051
rect 110029 239023 110064 239051
rect 109904 238989 110064 239023
rect 109904 238961 109939 238989
rect 109967 238961 110001 238989
rect 110029 238961 110064 238989
rect 109904 238944 110064 238961
rect 125264 239175 125424 239192
rect 125264 239147 125299 239175
rect 125327 239147 125361 239175
rect 125389 239147 125424 239175
rect 125264 239113 125424 239147
rect 125264 239085 125299 239113
rect 125327 239085 125361 239113
rect 125389 239085 125424 239113
rect 125264 239051 125424 239085
rect 125264 239023 125299 239051
rect 125327 239023 125361 239051
rect 125389 239023 125424 239051
rect 125264 238989 125424 239023
rect 125264 238961 125299 238989
rect 125327 238961 125361 238989
rect 125389 238961 125424 238989
rect 125264 238944 125424 238961
rect 140624 239175 140784 239192
rect 140624 239147 140659 239175
rect 140687 239147 140721 239175
rect 140749 239147 140784 239175
rect 140624 239113 140784 239147
rect 140624 239085 140659 239113
rect 140687 239085 140721 239113
rect 140749 239085 140784 239113
rect 140624 239051 140784 239085
rect 140624 239023 140659 239051
rect 140687 239023 140721 239051
rect 140749 239023 140784 239051
rect 140624 238989 140784 239023
rect 140624 238961 140659 238989
rect 140687 238961 140721 238989
rect 140749 238961 140784 238989
rect 140624 238944 140784 238961
rect 155984 239175 156144 239192
rect 155984 239147 156019 239175
rect 156047 239147 156081 239175
rect 156109 239147 156144 239175
rect 155984 239113 156144 239147
rect 155984 239085 156019 239113
rect 156047 239085 156081 239113
rect 156109 239085 156144 239113
rect 155984 239051 156144 239085
rect 155984 239023 156019 239051
rect 156047 239023 156081 239051
rect 156109 239023 156144 239051
rect 155984 238989 156144 239023
rect 155984 238961 156019 238989
rect 156047 238961 156081 238989
rect 156109 238961 156144 238989
rect 155984 238944 156144 238961
rect 102224 236175 102384 236192
rect 102224 236147 102259 236175
rect 102287 236147 102321 236175
rect 102349 236147 102384 236175
rect 102224 236113 102384 236147
rect 102224 236085 102259 236113
rect 102287 236085 102321 236113
rect 102349 236085 102384 236113
rect 102224 236051 102384 236085
rect 102224 236023 102259 236051
rect 102287 236023 102321 236051
rect 102349 236023 102384 236051
rect 102224 235989 102384 236023
rect 102224 235961 102259 235989
rect 102287 235961 102321 235989
rect 102349 235961 102384 235989
rect 102224 235944 102384 235961
rect 117584 236175 117744 236192
rect 117584 236147 117619 236175
rect 117647 236147 117681 236175
rect 117709 236147 117744 236175
rect 117584 236113 117744 236147
rect 117584 236085 117619 236113
rect 117647 236085 117681 236113
rect 117709 236085 117744 236113
rect 117584 236051 117744 236085
rect 117584 236023 117619 236051
rect 117647 236023 117681 236051
rect 117709 236023 117744 236051
rect 117584 235989 117744 236023
rect 117584 235961 117619 235989
rect 117647 235961 117681 235989
rect 117709 235961 117744 235989
rect 117584 235944 117744 235961
rect 132944 236175 133104 236192
rect 132944 236147 132979 236175
rect 133007 236147 133041 236175
rect 133069 236147 133104 236175
rect 132944 236113 133104 236147
rect 132944 236085 132979 236113
rect 133007 236085 133041 236113
rect 133069 236085 133104 236113
rect 132944 236051 133104 236085
rect 132944 236023 132979 236051
rect 133007 236023 133041 236051
rect 133069 236023 133104 236051
rect 132944 235989 133104 236023
rect 132944 235961 132979 235989
rect 133007 235961 133041 235989
rect 133069 235961 133104 235989
rect 132944 235944 133104 235961
rect 148304 236175 148464 236192
rect 148304 236147 148339 236175
rect 148367 236147 148401 236175
rect 148429 236147 148464 236175
rect 148304 236113 148464 236147
rect 148304 236085 148339 236113
rect 148367 236085 148401 236113
rect 148429 236085 148464 236113
rect 148304 236051 148464 236085
rect 148304 236023 148339 236051
rect 148367 236023 148401 236051
rect 148429 236023 148464 236051
rect 148304 235989 148464 236023
rect 148304 235961 148339 235989
rect 148367 235961 148401 235989
rect 148429 235961 148464 235989
rect 148304 235944 148464 235961
rect 163664 236175 163824 236192
rect 163664 236147 163699 236175
rect 163727 236147 163761 236175
rect 163789 236147 163824 236175
rect 163664 236113 163824 236147
rect 163664 236085 163699 236113
rect 163727 236085 163761 236113
rect 163789 236085 163824 236113
rect 163664 236051 163824 236085
rect 163664 236023 163699 236051
rect 163727 236023 163761 236051
rect 163789 236023 163824 236051
rect 163664 235989 163824 236023
rect 163664 235961 163699 235989
rect 163727 235961 163761 235989
rect 163789 235961 163824 235989
rect 163664 235944 163824 235961
rect 171669 236175 171979 244961
rect 171669 236147 171717 236175
rect 171745 236147 171779 236175
rect 171807 236147 171841 236175
rect 171869 236147 171903 236175
rect 171931 236147 171979 236175
rect 171669 236113 171979 236147
rect 171669 236085 171717 236113
rect 171745 236085 171779 236113
rect 171807 236085 171841 236113
rect 171869 236085 171903 236113
rect 171931 236085 171979 236113
rect 171669 236051 171979 236085
rect 171669 236023 171717 236051
rect 171745 236023 171779 236051
rect 171807 236023 171841 236051
rect 171869 236023 171903 236051
rect 171931 236023 171979 236051
rect 171669 235989 171979 236023
rect 171669 235961 171717 235989
rect 171745 235961 171779 235989
rect 171807 235961 171841 235989
rect 171869 235961 171903 235989
rect 171931 235961 171979 235989
rect 96729 230147 96777 230175
rect 96805 230147 96839 230175
rect 96867 230147 96901 230175
rect 96929 230147 96963 230175
rect 96991 230147 97039 230175
rect 96729 230113 97039 230147
rect 96729 230085 96777 230113
rect 96805 230085 96839 230113
rect 96867 230085 96901 230113
rect 96929 230085 96963 230113
rect 96991 230085 97039 230113
rect 96729 230051 97039 230085
rect 96729 230023 96777 230051
rect 96805 230023 96839 230051
rect 96867 230023 96901 230051
rect 96929 230023 96963 230051
rect 96991 230023 97039 230051
rect 96729 229989 97039 230023
rect 96729 229961 96777 229989
rect 96805 229961 96839 229989
rect 96867 229961 96901 229989
rect 96929 229961 96963 229989
rect 96991 229961 97039 229989
rect 96729 221175 97039 229961
rect 109904 230175 110064 230192
rect 109904 230147 109939 230175
rect 109967 230147 110001 230175
rect 110029 230147 110064 230175
rect 109904 230113 110064 230147
rect 109904 230085 109939 230113
rect 109967 230085 110001 230113
rect 110029 230085 110064 230113
rect 109904 230051 110064 230085
rect 109904 230023 109939 230051
rect 109967 230023 110001 230051
rect 110029 230023 110064 230051
rect 109904 229989 110064 230023
rect 109904 229961 109939 229989
rect 109967 229961 110001 229989
rect 110029 229961 110064 229989
rect 109904 229944 110064 229961
rect 125264 230175 125424 230192
rect 125264 230147 125299 230175
rect 125327 230147 125361 230175
rect 125389 230147 125424 230175
rect 125264 230113 125424 230147
rect 125264 230085 125299 230113
rect 125327 230085 125361 230113
rect 125389 230085 125424 230113
rect 125264 230051 125424 230085
rect 125264 230023 125299 230051
rect 125327 230023 125361 230051
rect 125389 230023 125424 230051
rect 125264 229989 125424 230023
rect 125264 229961 125299 229989
rect 125327 229961 125361 229989
rect 125389 229961 125424 229989
rect 125264 229944 125424 229961
rect 140624 230175 140784 230192
rect 140624 230147 140659 230175
rect 140687 230147 140721 230175
rect 140749 230147 140784 230175
rect 140624 230113 140784 230147
rect 140624 230085 140659 230113
rect 140687 230085 140721 230113
rect 140749 230085 140784 230113
rect 140624 230051 140784 230085
rect 140624 230023 140659 230051
rect 140687 230023 140721 230051
rect 140749 230023 140784 230051
rect 140624 229989 140784 230023
rect 140624 229961 140659 229989
rect 140687 229961 140721 229989
rect 140749 229961 140784 229989
rect 140624 229944 140784 229961
rect 155984 230175 156144 230192
rect 155984 230147 156019 230175
rect 156047 230147 156081 230175
rect 156109 230147 156144 230175
rect 155984 230113 156144 230147
rect 155984 230085 156019 230113
rect 156047 230085 156081 230113
rect 156109 230085 156144 230113
rect 155984 230051 156144 230085
rect 155984 230023 156019 230051
rect 156047 230023 156081 230051
rect 156109 230023 156144 230051
rect 155984 229989 156144 230023
rect 155984 229961 156019 229989
rect 156047 229961 156081 229989
rect 156109 229961 156144 229989
rect 155984 229944 156144 229961
rect 102224 227175 102384 227192
rect 102224 227147 102259 227175
rect 102287 227147 102321 227175
rect 102349 227147 102384 227175
rect 102224 227113 102384 227147
rect 102224 227085 102259 227113
rect 102287 227085 102321 227113
rect 102349 227085 102384 227113
rect 102224 227051 102384 227085
rect 102224 227023 102259 227051
rect 102287 227023 102321 227051
rect 102349 227023 102384 227051
rect 102224 226989 102384 227023
rect 102224 226961 102259 226989
rect 102287 226961 102321 226989
rect 102349 226961 102384 226989
rect 102224 226944 102384 226961
rect 117584 227175 117744 227192
rect 117584 227147 117619 227175
rect 117647 227147 117681 227175
rect 117709 227147 117744 227175
rect 117584 227113 117744 227147
rect 117584 227085 117619 227113
rect 117647 227085 117681 227113
rect 117709 227085 117744 227113
rect 117584 227051 117744 227085
rect 117584 227023 117619 227051
rect 117647 227023 117681 227051
rect 117709 227023 117744 227051
rect 117584 226989 117744 227023
rect 117584 226961 117619 226989
rect 117647 226961 117681 226989
rect 117709 226961 117744 226989
rect 117584 226944 117744 226961
rect 132944 227175 133104 227192
rect 132944 227147 132979 227175
rect 133007 227147 133041 227175
rect 133069 227147 133104 227175
rect 132944 227113 133104 227147
rect 132944 227085 132979 227113
rect 133007 227085 133041 227113
rect 133069 227085 133104 227113
rect 132944 227051 133104 227085
rect 132944 227023 132979 227051
rect 133007 227023 133041 227051
rect 133069 227023 133104 227051
rect 132944 226989 133104 227023
rect 132944 226961 132979 226989
rect 133007 226961 133041 226989
rect 133069 226961 133104 226989
rect 132944 226944 133104 226961
rect 148304 227175 148464 227192
rect 148304 227147 148339 227175
rect 148367 227147 148401 227175
rect 148429 227147 148464 227175
rect 148304 227113 148464 227147
rect 148304 227085 148339 227113
rect 148367 227085 148401 227113
rect 148429 227085 148464 227113
rect 148304 227051 148464 227085
rect 148304 227023 148339 227051
rect 148367 227023 148401 227051
rect 148429 227023 148464 227051
rect 148304 226989 148464 227023
rect 148304 226961 148339 226989
rect 148367 226961 148401 226989
rect 148429 226961 148464 226989
rect 148304 226944 148464 226961
rect 163664 227175 163824 227192
rect 163664 227147 163699 227175
rect 163727 227147 163761 227175
rect 163789 227147 163824 227175
rect 163664 227113 163824 227147
rect 163664 227085 163699 227113
rect 163727 227085 163761 227113
rect 163789 227085 163824 227113
rect 163664 227051 163824 227085
rect 163664 227023 163699 227051
rect 163727 227023 163761 227051
rect 163789 227023 163824 227051
rect 163664 226989 163824 227023
rect 163664 226961 163699 226989
rect 163727 226961 163761 226989
rect 163789 226961 163824 226989
rect 163664 226944 163824 226961
rect 171669 227175 171979 235961
rect 171669 227147 171717 227175
rect 171745 227147 171779 227175
rect 171807 227147 171841 227175
rect 171869 227147 171903 227175
rect 171931 227147 171979 227175
rect 171669 227113 171979 227147
rect 171669 227085 171717 227113
rect 171745 227085 171779 227113
rect 171807 227085 171841 227113
rect 171869 227085 171903 227113
rect 171931 227085 171979 227113
rect 171669 227051 171979 227085
rect 171669 227023 171717 227051
rect 171745 227023 171779 227051
rect 171807 227023 171841 227051
rect 171869 227023 171903 227051
rect 171931 227023 171979 227051
rect 171669 226989 171979 227023
rect 171669 226961 171717 226989
rect 171745 226961 171779 226989
rect 171807 226961 171841 226989
rect 171869 226961 171903 226989
rect 171931 226961 171979 226989
rect 96729 221147 96777 221175
rect 96805 221147 96839 221175
rect 96867 221147 96901 221175
rect 96929 221147 96963 221175
rect 96991 221147 97039 221175
rect 96729 221113 97039 221147
rect 96729 221085 96777 221113
rect 96805 221085 96839 221113
rect 96867 221085 96901 221113
rect 96929 221085 96963 221113
rect 96991 221085 97039 221113
rect 96729 221051 97039 221085
rect 96729 221023 96777 221051
rect 96805 221023 96839 221051
rect 96867 221023 96901 221051
rect 96929 221023 96963 221051
rect 96991 221023 97039 221051
rect 96729 220989 97039 221023
rect 96729 220961 96777 220989
rect 96805 220961 96839 220989
rect 96867 220961 96901 220989
rect 96929 220961 96963 220989
rect 96991 220961 97039 220989
rect 96729 212175 97039 220961
rect 109904 221175 110064 221192
rect 109904 221147 109939 221175
rect 109967 221147 110001 221175
rect 110029 221147 110064 221175
rect 109904 221113 110064 221147
rect 109904 221085 109939 221113
rect 109967 221085 110001 221113
rect 110029 221085 110064 221113
rect 109904 221051 110064 221085
rect 109904 221023 109939 221051
rect 109967 221023 110001 221051
rect 110029 221023 110064 221051
rect 109904 220989 110064 221023
rect 109904 220961 109939 220989
rect 109967 220961 110001 220989
rect 110029 220961 110064 220989
rect 109904 220944 110064 220961
rect 125264 221175 125424 221192
rect 125264 221147 125299 221175
rect 125327 221147 125361 221175
rect 125389 221147 125424 221175
rect 125264 221113 125424 221147
rect 125264 221085 125299 221113
rect 125327 221085 125361 221113
rect 125389 221085 125424 221113
rect 125264 221051 125424 221085
rect 125264 221023 125299 221051
rect 125327 221023 125361 221051
rect 125389 221023 125424 221051
rect 125264 220989 125424 221023
rect 125264 220961 125299 220989
rect 125327 220961 125361 220989
rect 125389 220961 125424 220989
rect 125264 220944 125424 220961
rect 140624 221175 140784 221192
rect 140624 221147 140659 221175
rect 140687 221147 140721 221175
rect 140749 221147 140784 221175
rect 140624 221113 140784 221147
rect 140624 221085 140659 221113
rect 140687 221085 140721 221113
rect 140749 221085 140784 221113
rect 140624 221051 140784 221085
rect 140624 221023 140659 221051
rect 140687 221023 140721 221051
rect 140749 221023 140784 221051
rect 140624 220989 140784 221023
rect 140624 220961 140659 220989
rect 140687 220961 140721 220989
rect 140749 220961 140784 220989
rect 140624 220944 140784 220961
rect 155984 221175 156144 221192
rect 155984 221147 156019 221175
rect 156047 221147 156081 221175
rect 156109 221147 156144 221175
rect 155984 221113 156144 221147
rect 155984 221085 156019 221113
rect 156047 221085 156081 221113
rect 156109 221085 156144 221113
rect 155984 221051 156144 221085
rect 155984 221023 156019 221051
rect 156047 221023 156081 221051
rect 156109 221023 156144 221051
rect 155984 220989 156144 221023
rect 155984 220961 156019 220989
rect 156047 220961 156081 220989
rect 156109 220961 156144 220989
rect 155984 220944 156144 220961
rect 102224 218175 102384 218192
rect 102224 218147 102259 218175
rect 102287 218147 102321 218175
rect 102349 218147 102384 218175
rect 102224 218113 102384 218147
rect 102224 218085 102259 218113
rect 102287 218085 102321 218113
rect 102349 218085 102384 218113
rect 102224 218051 102384 218085
rect 102224 218023 102259 218051
rect 102287 218023 102321 218051
rect 102349 218023 102384 218051
rect 102224 217989 102384 218023
rect 102224 217961 102259 217989
rect 102287 217961 102321 217989
rect 102349 217961 102384 217989
rect 102224 217944 102384 217961
rect 117584 218175 117744 218192
rect 117584 218147 117619 218175
rect 117647 218147 117681 218175
rect 117709 218147 117744 218175
rect 117584 218113 117744 218147
rect 117584 218085 117619 218113
rect 117647 218085 117681 218113
rect 117709 218085 117744 218113
rect 117584 218051 117744 218085
rect 117584 218023 117619 218051
rect 117647 218023 117681 218051
rect 117709 218023 117744 218051
rect 117584 217989 117744 218023
rect 117584 217961 117619 217989
rect 117647 217961 117681 217989
rect 117709 217961 117744 217989
rect 117584 217944 117744 217961
rect 132944 218175 133104 218192
rect 132944 218147 132979 218175
rect 133007 218147 133041 218175
rect 133069 218147 133104 218175
rect 132944 218113 133104 218147
rect 132944 218085 132979 218113
rect 133007 218085 133041 218113
rect 133069 218085 133104 218113
rect 132944 218051 133104 218085
rect 132944 218023 132979 218051
rect 133007 218023 133041 218051
rect 133069 218023 133104 218051
rect 132944 217989 133104 218023
rect 132944 217961 132979 217989
rect 133007 217961 133041 217989
rect 133069 217961 133104 217989
rect 132944 217944 133104 217961
rect 148304 218175 148464 218192
rect 148304 218147 148339 218175
rect 148367 218147 148401 218175
rect 148429 218147 148464 218175
rect 148304 218113 148464 218147
rect 148304 218085 148339 218113
rect 148367 218085 148401 218113
rect 148429 218085 148464 218113
rect 148304 218051 148464 218085
rect 148304 218023 148339 218051
rect 148367 218023 148401 218051
rect 148429 218023 148464 218051
rect 148304 217989 148464 218023
rect 148304 217961 148339 217989
rect 148367 217961 148401 217989
rect 148429 217961 148464 217989
rect 148304 217944 148464 217961
rect 163664 218175 163824 218192
rect 163664 218147 163699 218175
rect 163727 218147 163761 218175
rect 163789 218147 163824 218175
rect 163664 218113 163824 218147
rect 163664 218085 163699 218113
rect 163727 218085 163761 218113
rect 163789 218085 163824 218113
rect 163664 218051 163824 218085
rect 163664 218023 163699 218051
rect 163727 218023 163761 218051
rect 163789 218023 163824 218051
rect 163664 217989 163824 218023
rect 163664 217961 163699 217989
rect 163727 217961 163761 217989
rect 163789 217961 163824 217989
rect 163664 217944 163824 217961
rect 171669 218175 171979 226961
rect 171669 218147 171717 218175
rect 171745 218147 171779 218175
rect 171807 218147 171841 218175
rect 171869 218147 171903 218175
rect 171931 218147 171979 218175
rect 171669 218113 171979 218147
rect 171669 218085 171717 218113
rect 171745 218085 171779 218113
rect 171807 218085 171841 218113
rect 171869 218085 171903 218113
rect 171931 218085 171979 218113
rect 171669 218051 171979 218085
rect 171669 218023 171717 218051
rect 171745 218023 171779 218051
rect 171807 218023 171841 218051
rect 171869 218023 171903 218051
rect 171931 218023 171979 218051
rect 171669 217989 171979 218023
rect 171669 217961 171717 217989
rect 171745 217961 171779 217989
rect 171807 217961 171841 217989
rect 171869 217961 171903 217989
rect 171931 217961 171979 217989
rect 96729 212147 96777 212175
rect 96805 212147 96839 212175
rect 96867 212147 96901 212175
rect 96929 212147 96963 212175
rect 96991 212147 97039 212175
rect 96729 212113 97039 212147
rect 96729 212085 96777 212113
rect 96805 212085 96839 212113
rect 96867 212085 96901 212113
rect 96929 212085 96963 212113
rect 96991 212085 97039 212113
rect 96729 212051 97039 212085
rect 96729 212023 96777 212051
rect 96805 212023 96839 212051
rect 96867 212023 96901 212051
rect 96929 212023 96963 212051
rect 96991 212023 97039 212051
rect 96729 211989 97039 212023
rect 96729 211961 96777 211989
rect 96805 211961 96839 211989
rect 96867 211961 96901 211989
rect 96929 211961 96963 211989
rect 96991 211961 97039 211989
rect 96729 203175 97039 211961
rect 109904 212175 110064 212192
rect 109904 212147 109939 212175
rect 109967 212147 110001 212175
rect 110029 212147 110064 212175
rect 109904 212113 110064 212147
rect 109904 212085 109939 212113
rect 109967 212085 110001 212113
rect 110029 212085 110064 212113
rect 109904 212051 110064 212085
rect 109904 212023 109939 212051
rect 109967 212023 110001 212051
rect 110029 212023 110064 212051
rect 109904 211989 110064 212023
rect 109904 211961 109939 211989
rect 109967 211961 110001 211989
rect 110029 211961 110064 211989
rect 109904 211944 110064 211961
rect 125264 212175 125424 212192
rect 125264 212147 125299 212175
rect 125327 212147 125361 212175
rect 125389 212147 125424 212175
rect 125264 212113 125424 212147
rect 125264 212085 125299 212113
rect 125327 212085 125361 212113
rect 125389 212085 125424 212113
rect 125264 212051 125424 212085
rect 125264 212023 125299 212051
rect 125327 212023 125361 212051
rect 125389 212023 125424 212051
rect 125264 211989 125424 212023
rect 125264 211961 125299 211989
rect 125327 211961 125361 211989
rect 125389 211961 125424 211989
rect 125264 211944 125424 211961
rect 140624 212175 140784 212192
rect 140624 212147 140659 212175
rect 140687 212147 140721 212175
rect 140749 212147 140784 212175
rect 140624 212113 140784 212147
rect 140624 212085 140659 212113
rect 140687 212085 140721 212113
rect 140749 212085 140784 212113
rect 140624 212051 140784 212085
rect 140624 212023 140659 212051
rect 140687 212023 140721 212051
rect 140749 212023 140784 212051
rect 140624 211989 140784 212023
rect 140624 211961 140659 211989
rect 140687 211961 140721 211989
rect 140749 211961 140784 211989
rect 140624 211944 140784 211961
rect 155984 212175 156144 212192
rect 155984 212147 156019 212175
rect 156047 212147 156081 212175
rect 156109 212147 156144 212175
rect 155984 212113 156144 212147
rect 155984 212085 156019 212113
rect 156047 212085 156081 212113
rect 156109 212085 156144 212113
rect 155984 212051 156144 212085
rect 155984 212023 156019 212051
rect 156047 212023 156081 212051
rect 156109 212023 156144 212051
rect 155984 211989 156144 212023
rect 155984 211961 156019 211989
rect 156047 211961 156081 211989
rect 156109 211961 156144 211989
rect 155984 211944 156144 211961
rect 102224 209175 102384 209192
rect 102224 209147 102259 209175
rect 102287 209147 102321 209175
rect 102349 209147 102384 209175
rect 102224 209113 102384 209147
rect 102224 209085 102259 209113
rect 102287 209085 102321 209113
rect 102349 209085 102384 209113
rect 102224 209051 102384 209085
rect 102224 209023 102259 209051
rect 102287 209023 102321 209051
rect 102349 209023 102384 209051
rect 102224 208989 102384 209023
rect 102224 208961 102259 208989
rect 102287 208961 102321 208989
rect 102349 208961 102384 208989
rect 102224 208944 102384 208961
rect 117584 209175 117744 209192
rect 117584 209147 117619 209175
rect 117647 209147 117681 209175
rect 117709 209147 117744 209175
rect 117584 209113 117744 209147
rect 117584 209085 117619 209113
rect 117647 209085 117681 209113
rect 117709 209085 117744 209113
rect 117584 209051 117744 209085
rect 117584 209023 117619 209051
rect 117647 209023 117681 209051
rect 117709 209023 117744 209051
rect 117584 208989 117744 209023
rect 117584 208961 117619 208989
rect 117647 208961 117681 208989
rect 117709 208961 117744 208989
rect 117584 208944 117744 208961
rect 132944 209175 133104 209192
rect 132944 209147 132979 209175
rect 133007 209147 133041 209175
rect 133069 209147 133104 209175
rect 132944 209113 133104 209147
rect 132944 209085 132979 209113
rect 133007 209085 133041 209113
rect 133069 209085 133104 209113
rect 132944 209051 133104 209085
rect 132944 209023 132979 209051
rect 133007 209023 133041 209051
rect 133069 209023 133104 209051
rect 132944 208989 133104 209023
rect 132944 208961 132979 208989
rect 133007 208961 133041 208989
rect 133069 208961 133104 208989
rect 132944 208944 133104 208961
rect 148304 209175 148464 209192
rect 148304 209147 148339 209175
rect 148367 209147 148401 209175
rect 148429 209147 148464 209175
rect 148304 209113 148464 209147
rect 148304 209085 148339 209113
rect 148367 209085 148401 209113
rect 148429 209085 148464 209113
rect 148304 209051 148464 209085
rect 148304 209023 148339 209051
rect 148367 209023 148401 209051
rect 148429 209023 148464 209051
rect 148304 208989 148464 209023
rect 148304 208961 148339 208989
rect 148367 208961 148401 208989
rect 148429 208961 148464 208989
rect 148304 208944 148464 208961
rect 163664 209175 163824 209192
rect 163664 209147 163699 209175
rect 163727 209147 163761 209175
rect 163789 209147 163824 209175
rect 163664 209113 163824 209147
rect 163664 209085 163699 209113
rect 163727 209085 163761 209113
rect 163789 209085 163824 209113
rect 163664 209051 163824 209085
rect 163664 209023 163699 209051
rect 163727 209023 163761 209051
rect 163789 209023 163824 209051
rect 163664 208989 163824 209023
rect 163664 208961 163699 208989
rect 163727 208961 163761 208989
rect 163789 208961 163824 208989
rect 163664 208944 163824 208961
rect 171669 209175 171979 217961
rect 171669 209147 171717 209175
rect 171745 209147 171779 209175
rect 171807 209147 171841 209175
rect 171869 209147 171903 209175
rect 171931 209147 171979 209175
rect 171669 209113 171979 209147
rect 171669 209085 171717 209113
rect 171745 209085 171779 209113
rect 171807 209085 171841 209113
rect 171869 209085 171903 209113
rect 171931 209085 171979 209113
rect 171669 209051 171979 209085
rect 171669 209023 171717 209051
rect 171745 209023 171779 209051
rect 171807 209023 171841 209051
rect 171869 209023 171903 209051
rect 171931 209023 171979 209051
rect 171669 208989 171979 209023
rect 171669 208961 171717 208989
rect 171745 208961 171779 208989
rect 171807 208961 171841 208989
rect 171869 208961 171903 208989
rect 171931 208961 171979 208989
rect 96729 203147 96777 203175
rect 96805 203147 96839 203175
rect 96867 203147 96901 203175
rect 96929 203147 96963 203175
rect 96991 203147 97039 203175
rect 96729 203113 97039 203147
rect 96729 203085 96777 203113
rect 96805 203085 96839 203113
rect 96867 203085 96901 203113
rect 96929 203085 96963 203113
rect 96991 203085 97039 203113
rect 96729 203051 97039 203085
rect 96729 203023 96777 203051
rect 96805 203023 96839 203051
rect 96867 203023 96901 203051
rect 96929 203023 96963 203051
rect 96991 203023 97039 203051
rect 96729 202989 97039 203023
rect 96729 202961 96777 202989
rect 96805 202961 96839 202989
rect 96867 202961 96901 202989
rect 96929 202961 96963 202989
rect 96991 202961 97039 202989
rect 96729 194175 97039 202961
rect 109904 203175 110064 203192
rect 109904 203147 109939 203175
rect 109967 203147 110001 203175
rect 110029 203147 110064 203175
rect 109904 203113 110064 203147
rect 109904 203085 109939 203113
rect 109967 203085 110001 203113
rect 110029 203085 110064 203113
rect 109904 203051 110064 203085
rect 109904 203023 109939 203051
rect 109967 203023 110001 203051
rect 110029 203023 110064 203051
rect 109904 202989 110064 203023
rect 109904 202961 109939 202989
rect 109967 202961 110001 202989
rect 110029 202961 110064 202989
rect 109904 202944 110064 202961
rect 125264 203175 125424 203192
rect 125264 203147 125299 203175
rect 125327 203147 125361 203175
rect 125389 203147 125424 203175
rect 125264 203113 125424 203147
rect 125264 203085 125299 203113
rect 125327 203085 125361 203113
rect 125389 203085 125424 203113
rect 125264 203051 125424 203085
rect 125264 203023 125299 203051
rect 125327 203023 125361 203051
rect 125389 203023 125424 203051
rect 125264 202989 125424 203023
rect 125264 202961 125299 202989
rect 125327 202961 125361 202989
rect 125389 202961 125424 202989
rect 125264 202944 125424 202961
rect 140624 203175 140784 203192
rect 140624 203147 140659 203175
rect 140687 203147 140721 203175
rect 140749 203147 140784 203175
rect 140624 203113 140784 203147
rect 140624 203085 140659 203113
rect 140687 203085 140721 203113
rect 140749 203085 140784 203113
rect 140624 203051 140784 203085
rect 140624 203023 140659 203051
rect 140687 203023 140721 203051
rect 140749 203023 140784 203051
rect 140624 202989 140784 203023
rect 140624 202961 140659 202989
rect 140687 202961 140721 202989
rect 140749 202961 140784 202989
rect 140624 202944 140784 202961
rect 155984 203175 156144 203192
rect 155984 203147 156019 203175
rect 156047 203147 156081 203175
rect 156109 203147 156144 203175
rect 155984 203113 156144 203147
rect 155984 203085 156019 203113
rect 156047 203085 156081 203113
rect 156109 203085 156144 203113
rect 155984 203051 156144 203085
rect 155984 203023 156019 203051
rect 156047 203023 156081 203051
rect 156109 203023 156144 203051
rect 155984 202989 156144 203023
rect 155984 202961 156019 202989
rect 156047 202961 156081 202989
rect 156109 202961 156144 202989
rect 155984 202944 156144 202961
rect 102224 200175 102384 200192
rect 102224 200147 102259 200175
rect 102287 200147 102321 200175
rect 102349 200147 102384 200175
rect 102224 200113 102384 200147
rect 102224 200085 102259 200113
rect 102287 200085 102321 200113
rect 102349 200085 102384 200113
rect 102224 200051 102384 200085
rect 102224 200023 102259 200051
rect 102287 200023 102321 200051
rect 102349 200023 102384 200051
rect 102224 199989 102384 200023
rect 102224 199961 102259 199989
rect 102287 199961 102321 199989
rect 102349 199961 102384 199989
rect 102224 199944 102384 199961
rect 117584 200175 117744 200192
rect 117584 200147 117619 200175
rect 117647 200147 117681 200175
rect 117709 200147 117744 200175
rect 117584 200113 117744 200147
rect 117584 200085 117619 200113
rect 117647 200085 117681 200113
rect 117709 200085 117744 200113
rect 117584 200051 117744 200085
rect 117584 200023 117619 200051
rect 117647 200023 117681 200051
rect 117709 200023 117744 200051
rect 117584 199989 117744 200023
rect 117584 199961 117619 199989
rect 117647 199961 117681 199989
rect 117709 199961 117744 199989
rect 117584 199944 117744 199961
rect 132944 200175 133104 200192
rect 132944 200147 132979 200175
rect 133007 200147 133041 200175
rect 133069 200147 133104 200175
rect 132944 200113 133104 200147
rect 132944 200085 132979 200113
rect 133007 200085 133041 200113
rect 133069 200085 133104 200113
rect 132944 200051 133104 200085
rect 132944 200023 132979 200051
rect 133007 200023 133041 200051
rect 133069 200023 133104 200051
rect 132944 199989 133104 200023
rect 132944 199961 132979 199989
rect 133007 199961 133041 199989
rect 133069 199961 133104 199989
rect 132944 199944 133104 199961
rect 148304 200175 148464 200192
rect 148304 200147 148339 200175
rect 148367 200147 148401 200175
rect 148429 200147 148464 200175
rect 148304 200113 148464 200147
rect 148304 200085 148339 200113
rect 148367 200085 148401 200113
rect 148429 200085 148464 200113
rect 148304 200051 148464 200085
rect 148304 200023 148339 200051
rect 148367 200023 148401 200051
rect 148429 200023 148464 200051
rect 148304 199989 148464 200023
rect 148304 199961 148339 199989
rect 148367 199961 148401 199989
rect 148429 199961 148464 199989
rect 148304 199944 148464 199961
rect 163664 200175 163824 200192
rect 163664 200147 163699 200175
rect 163727 200147 163761 200175
rect 163789 200147 163824 200175
rect 163664 200113 163824 200147
rect 163664 200085 163699 200113
rect 163727 200085 163761 200113
rect 163789 200085 163824 200113
rect 163664 200051 163824 200085
rect 163664 200023 163699 200051
rect 163727 200023 163761 200051
rect 163789 200023 163824 200051
rect 163664 199989 163824 200023
rect 163664 199961 163699 199989
rect 163727 199961 163761 199989
rect 163789 199961 163824 199989
rect 163664 199944 163824 199961
rect 171669 200175 171979 208961
rect 171669 200147 171717 200175
rect 171745 200147 171779 200175
rect 171807 200147 171841 200175
rect 171869 200147 171903 200175
rect 171931 200147 171979 200175
rect 171669 200113 171979 200147
rect 171669 200085 171717 200113
rect 171745 200085 171779 200113
rect 171807 200085 171841 200113
rect 171869 200085 171903 200113
rect 171931 200085 171979 200113
rect 171669 200051 171979 200085
rect 171669 200023 171717 200051
rect 171745 200023 171779 200051
rect 171807 200023 171841 200051
rect 171869 200023 171903 200051
rect 171931 200023 171979 200051
rect 171669 199989 171979 200023
rect 171669 199961 171717 199989
rect 171745 199961 171779 199989
rect 171807 199961 171841 199989
rect 171869 199961 171903 199989
rect 171931 199961 171979 199989
rect 96729 194147 96777 194175
rect 96805 194147 96839 194175
rect 96867 194147 96901 194175
rect 96929 194147 96963 194175
rect 96991 194147 97039 194175
rect 96729 194113 97039 194147
rect 96729 194085 96777 194113
rect 96805 194085 96839 194113
rect 96867 194085 96901 194113
rect 96929 194085 96963 194113
rect 96991 194085 97039 194113
rect 96729 194051 97039 194085
rect 96729 194023 96777 194051
rect 96805 194023 96839 194051
rect 96867 194023 96901 194051
rect 96929 194023 96963 194051
rect 96991 194023 97039 194051
rect 96729 193989 97039 194023
rect 96729 193961 96777 193989
rect 96805 193961 96839 193989
rect 96867 193961 96901 193989
rect 96929 193961 96963 193989
rect 96991 193961 97039 193989
rect 96729 185175 97039 193961
rect 109904 194175 110064 194192
rect 109904 194147 109939 194175
rect 109967 194147 110001 194175
rect 110029 194147 110064 194175
rect 109904 194113 110064 194147
rect 109904 194085 109939 194113
rect 109967 194085 110001 194113
rect 110029 194085 110064 194113
rect 109904 194051 110064 194085
rect 109904 194023 109939 194051
rect 109967 194023 110001 194051
rect 110029 194023 110064 194051
rect 109904 193989 110064 194023
rect 109904 193961 109939 193989
rect 109967 193961 110001 193989
rect 110029 193961 110064 193989
rect 109904 193944 110064 193961
rect 125264 194175 125424 194192
rect 125264 194147 125299 194175
rect 125327 194147 125361 194175
rect 125389 194147 125424 194175
rect 125264 194113 125424 194147
rect 125264 194085 125299 194113
rect 125327 194085 125361 194113
rect 125389 194085 125424 194113
rect 125264 194051 125424 194085
rect 125264 194023 125299 194051
rect 125327 194023 125361 194051
rect 125389 194023 125424 194051
rect 125264 193989 125424 194023
rect 125264 193961 125299 193989
rect 125327 193961 125361 193989
rect 125389 193961 125424 193989
rect 125264 193944 125424 193961
rect 140624 194175 140784 194192
rect 140624 194147 140659 194175
rect 140687 194147 140721 194175
rect 140749 194147 140784 194175
rect 140624 194113 140784 194147
rect 140624 194085 140659 194113
rect 140687 194085 140721 194113
rect 140749 194085 140784 194113
rect 140624 194051 140784 194085
rect 140624 194023 140659 194051
rect 140687 194023 140721 194051
rect 140749 194023 140784 194051
rect 140624 193989 140784 194023
rect 140624 193961 140659 193989
rect 140687 193961 140721 193989
rect 140749 193961 140784 193989
rect 140624 193944 140784 193961
rect 155984 194175 156144 194192
rect 155984 194147 156019 194175
rect 156047 194147 156081 194175
rect 156109 194147 156144 194175
rect 155984 194113 156144 194147
rect 155984 194085 156019 194113
rect 156047 194085 156081 194113
rect 156109 194085 156144 194113
rect 155984 194051 156144 194085
rect 155984 194023 156019 194051
rect 156047 194023 156081 194051
rect 156109 194023 156144 194051
rect 155984 193989 156144 194023
rect 155984 193961 156019 193989
rect 156047 193961 156081 193989
rect 156109 193961 156144 193989
rect 155984 193944 156144 193961
rect 102224 191175 102384 191192
rect 102224 191147 102259 191175
rect 102287 191147 102321 191175
rect 102349 191147 102384 191175
rect 102224 191113 102384 191147
rect 102224 191085 102259 191113
rect 102287 191085 102321 191113
rect 102349 191085 102384 191113
rect 102224 191051 102384 191085
rect 102224 191023 102259 191051
rect 102287 191023 102321 191051
rect 102349 191023 102384 191051
rect 102224 190989 102384 191023
rect 102224 190961 102259 190989
rect 102287 190961 102321 190989
rect 102349 190961 102384 190989
rect 102224 190944 102384 190961
rect 117584 191175 117744 191192
rect 117584 191147 117619 191175
rect 117647 191147 117681 191175
rect 117709 191147 117744 191175
rect 117584 191113 117744 191147
rect 117584 191085 117619 191113
rect 117647 191085 117681 191113
rect 117709 191085 117744 191113
rect 117584 191051 117744 191085
rect 117584 191023 117619 191051
rect 117647 191023 117681 191051
rect 117709 191023 117744 191051
rect 117584 190989 117744 191023
rect 117584 190961 117619 190989
rect 117647 190961 117681 190989
rect 117709 190961 117744 190989
rect 117584 190944 117744 190961
rect 132944 191175 133104 191192
rect 132944 191147 132979 191175
rect 133007 191147 133041 191175
rect 133069 191147 133104 191175
rect 132944 191113 133104 191147
rect 132944 191085 132979 191113
rect 133007 191085 133041 191113
rect 133069 191085 133104 191113
rect 132944 191051 133104 191085
rect 132944 191023 132979 191051
rect 133007 191023 133041 191051
rect 133069 191023 133104 191051
rect 132944 190989 133104 191023
rect 132944 190961 132979 190989
rect 133007 190961 133041 190989
rect 133069 190961 133104 190989
rect 132944 190944 133104 190961
rect 148304 191175 148464 191192
rect 148304 191147 148339 191175
rect 148367 191147 148401 191175
rect 148429 191147 148464 191175
rect 148304 191113 148464 191147
rect 148304 191085 148339 191113
rect 148367 191085 148401 191113
rect 148429 191085 148464 191113
rect 148304 191051 148464 191085
rect 148304 191023 148339 191051
rect 148367 191023 148401 191051
rect 148429 191023 148464 191051
rect 148304 190989 148464 191023
rect 148304 190961 148339 190989
rect 148367 190961 148401 190989
rect 148429 190961 148464 190989
rect 148304 190944 148464 190961
rect 163664 191175 163824 191192
rect 163664 191147 163699 191175
rect 163727 191147 163761 191175
rect 163789 191147 163824 191175
rect 163664 191113 163824 191147
rect 163664 191085 163699 191113
rect 163727 191085 163761 191113
rect 163789 191085 163824 191113
rect 163664 191051 163824 191085
rect 163664 191023 163699 191051
rect 163727 191023 163761 191051
rect 163789 191023 163824 191051
rect 163664 190989 163824 191023
rect 163664 190961 163699 190989
rect 163727 190961 163761 190989
rect 163789 190961 163824 190989
rect 163664 190944 163824 190961
rect 171669 191175 171979 199961
rect 171669 191147 171717 191175
rect 171745 191147 171779 191175
rect 171807 191147 171841 191175
rect 171869 191147 171903 191175
rect 171931 191147 171979 191175
rect 171669 191113 171979 191147
rect 171669 191085 171717 191113
rect 171745 191085 171779 191113
rect 171807 191085 171841 191113
rect 171869 191085 171903 191113
rect 171931 191085 171979 191113
rect 171669 191051 171979 191085
rect 171669 191023 171717 191051
rect 171745 191023 171779 191051
rect 171807 191023 171841 191051
rect 171869 191023 171903 191051
rect 171931 191023 171979 191051
rect 171669 190989 171979 191023
rect 171669 190961 171717 190989
rect 171745 190961 171779 190989
rect 171807 190961 171841 190989
rect 171869 190961 171903 190989
rect 171931 190961 171979 190989
rect 96729 185147 96777 185175
rect 96805 185147 96839 185175
rect 96867 185147 96901 185175
rect 96929 185147 96963 185175
rect 96991 185147 97039 185175
rect 96729 185113 97039 185147
rect 96729 185085 96777 185113
rect 96805 185085 96839 185113
rect 96867 185085 96901 185113
rect 96929 185085 96963 185113
rect 96991 185085 97039 185113
rect 96729 185051 97039 185085
rect 96729 185023 96777 185051
rect 96805 185023 96839 185051
rect 96867 185023 96901 185051
rect 96929 185023 96963 185051
rect 96991 185023 97039 185051
rect 96729 184989 97039 185023
rect 96729 184961 96777 184989
rect 96805 184961 96839 184989
rect 96867 184961 96901 184989
rect 96929 184961 96963 184989
rect 96991 184961 97039 184989
rect 96729 176175 97039 184961
rect 109904 185175 110064 185192
rect 109904 185147 109939 185175
rect 109967 185147 110001 185175
rect 110029 185147 110064 185175
rect 109904 185113 110064 185147
rect 109904 185085 109939 185113
rect 109967 185085 110001 185113
rect 110029 185085 110064 185113
rect 109904 185051 110064 185085
rect 109904 185023 109939 185051
rect 109967 185023 110001 185051
rect 110029 185023 110064 185051
rect 109904 184989 110064 185023
rect 109904 184961 109939 184989
rect 109967 184961 110001 184989
rect 110029 184961 110064 184989
rect 109904 184944 110064 184961
rect 125264 185175 125424 185192
rect 125264 185147 125299 185175
rect 125327 185147 125361 185175
rect 125389 185147 125424 185175
rect 125264 185113 125424 185147
rect 125264 185085 125299 185113
rect 125327 185085 125361 185113
rect 125389 185085 125424 185113
rect 125264 185051 125424 185085
rect 125264 185023 125299 185051
rect 125327 185023 125361 185051
rect 125389 185023 125424 185051
rect 125264 184989 125424 185023
rect 125264 184961 125299 184989
rect 125327 184961 125361 184989
rect 125389 184961 125424 184989
rect 125264 184944 125424 184961
rect 140624 185175 140784 185192
rect 140624 185147 140659 185175
rect 140687 185147 140721 185175
rect 140749 185147 140784 185175
rect 140624 185113 140784 185147
rect 140624 185085 140659 185113
rect 140687 185085 140721 185113
rect 140749 185085 140784 185113
rect 140624 185051 140784 185085
rect 140624 185023 140659 185051
rect 140687 185023 140721 185051
rect 140749 185023 140784 185051
rect 140624 184989 140784 185023
rect 140624 184961 140659 184989
rect 140687 184961 140721 184989
rect 140749 184961 140784 184989
rect 140624 184944 140784 184961
rect 155984 185175 156144 185192
rect 155984 185147 156019 185175
rect 156047 185147 156081 185175
rect 156109 185147 156144 185175
rect 155984 185113 156144 185147
rect 155984 185085 156019 185113
rect 156047 185085 156081 185113
rect 156109 185085 156144 185113
rect 155984 185051 156144 185085
rect 155984 185023 156019 185051
rect 156047 185023 156081 185051
rect 156109 185023 156144 185051
rect 155984 184989 156144 185023
rect 155984 184961 156019 184989
rect 156047 184961 156081 184989
rect 156109 184961 156144 184989
rect 155984 184944 156144 184961
rect 102224 182175 102384 182192
rect 102224 182147 102259 182175
rect 102287 182147 102321 182175
rect 102349 182147 102384 182175
rect 102224 182113 102384 182147
rect 102224 182085 102259 182113
rect 102287 182085 102321 182113
rect 102349 182085 102384 182113
rect 102224 182051 102384 182085
rect 102224 182023 102259 182051
rect 102287 182023 102321 182051
rect 102349 182023 102384 182051
rect 102224 181989 102384 182023
rect 102224 181961 102259 181989
rect 102287 181961 102321 181989
rect 102349 181961 102384 181989
rect 102224 181944 102384 181961
rect 117584 182175 117744 182192
rect 117584 182147 117619 182175
rect 117647 182147 117681 182175
rect 117709 182147 117744 182175
rect 117584 182113 117744 182147
rect 117584 182085 117619 182113
rect 117647 182085 117681 182113
rect 117709 182085 117744 182113
rect 117584 182051 117744 182085
rect 117584 182023 117619 182051
rect 117647 182023 117681 182051
rect 117709 182023 117744 182051
rect 117584 181989 117744 182023
rect 117584 181961 117619 181989
rect 117647 181961 117681 181989
rect 117709 181961 117744 181989
rect 117584 181944 117744 181961
rect 132944 182175 133104 182192
rect 132944 182147 132979 182175
rect 133007 182147 133041 182175
rect 133069 182147 133104 182175
rect 132944 182113 133104 182147
rect 132944 182085 132979 182113
rect 133007 182085 133041 182113
rect 133069 182085 133104 182113
rect 132944 182051 133104 182085
rect 132944 182023 132979 182051
rect 133007 182023 133041 182051
rect 133069 182023 133104 182051
rect 132944 181989 133104 182023
rect 132944 181961 132979 181989
rect 133007 181961 133041 181989
rect 133069 181961 133104 181989
rect 132944 181944 133104 181961
rect 148304 182175 148464 182192
rect 148304 182147 148339 182175
rect 148367 182147 148401 182175
rect 148429 182147 148464 182175
rect 148304 182113 148464 182147
rect 148304 182085 148339 182113
rect 148367 182085 148401 182113
rect 148429 182085 148464 182113
rect 148304 182051 148464 182085
rect 148304 182023 148339 182051
rect 148367 182023 148401 182051
rect 148429 182023 148464 182051
rect 148304 181989 148464 182023
rect 148304 181961 148339 181989
rect 148367 181961 148401 181989
rect 148429 181961 148464 181989
rect 148304 181944 148464 181961
rect 163664 182175 163824 182192
rect 163664 182147 163699 182175
rect 163727 182147 163761 182175
rect 163789 182147 163824 182175
rect 163664 182113 163824 182147
rect 163664 182085 163699 182113
rect 163727 182085 163761 182113
rect 163789 182085 163824 182113
rect 163664 182051 163824 182085
rect 163664 182023 163699 182051
rect 163727 182023 163761 182051
rect 163789 182023 163824 182051
rect 163664 181989 163824 182023
rect 163664 181961 163699 181989
rect 163727 181961 163761 181989
rect 163789 181961 163824 181989
rect 163664 181944 163824 181961
rect 171669 182175 171979 190961
rect 171669 182147 171717 182175
rect 171745 182147 171779 182175
rect 171807 182147 171841 182175
rect 171869 182147 171903 182175
rect 171931 182147 171979 182175
rect 171669 182113 171979 182147
rect 171669 182085 171717 182113
rect 171745 182085 171779 182113
rect 171807 182085 171841 182113
rect 171869 182085 171903 182113
rect 171931 182085 171979 182113
rect 171669 182051 171979 182085
rect 171669 182023 171717 182051
rect 171745 182023 171779 182051
rect 171807 182023 171841 182051
rect 171869 182023 171903 182051
rect 171931 182023 171979 182051
rect 171669 181989 171979 182023
rect 171669 181961 171717 181989
rect 171745 181961 171779 181989
rect 171807 181961 171841 181989
rect 171869 181961 171903 181989
rect 171931 181961 171979 181989
rect 96729 176147 96777 176175
rect 96805 176147 96839 176175
rect 96867 176147 96901 176175
rect 96929 176147 96963 176175
rect 96991 176147 97039 176175
rect 96729 176113 97039 176147
rect 96729 176085 96777 176113
rect 96805 176085 96839 176113
rect 96867 176085 96901 176113
rect 96929 176085 96963 176113
rect 96991 176085 97039 176113
rect 96729 176051 97039 176085
rect 96729 176023 96777 176051
rect 96805 176023 96839 176051
rect 96867 176023 96901 176051
rect 96929 176023 96963 176051
rect 96991 176023 97039 176051
rect 96729 175989 97039 176023
rect 96729 175961 96777 175989
rect 96805 175961 96839 175989
rect 96867 175961 96901 175989
rect 96929 175961 96963 175989
rect 96991 175961 97039 175989
rect 96729 167175 97039 175961
rect 109904 176175 110064 176192
rect 109904 176147 109939 176175
rect 109967 176147 110001 176175
rect 110029 176147 110064 176175
rect 109904 176113 110064 176147
rect 109904 176085 109939 176113
rect 109967 176085 110001 176113
rect 110029 176085 110064 176113
rect 109904 176051 110064 176085
rect 109904 176023 109939 176051
rect 109967 176023 110001 176051
rect 110029 176023 110064 176051
rect 109904 175989 110064 176023
rect 109904 175961 109939 175989
rect 109967 175961 110001 175989
rect 110029 175961 110064 175989
rect 109904 175944 110064 175961
rect 125264 176175 125424 176192
rect 125264 176147 125299 176175
rect 125327 176147 125361 176175
rect 125389 176147 125424 176175
rect 125264 176113 125424 176147
rect 125264 176085 125299 176113
rect 125327 176085 125361 176113
rect 125389 176085 125424 176113
rect 125264 176051 125424 176085
rect 125264 176023 125299 176051
rect 125327 176023 125361 176051
rect 125389 176023 125424 176051
rect 125264 175989 125424 176023
rect 125264 175961 125299 175989
rect 125327 175961 125361 175989
rect 125389 175961 125424 175989
rect 125264 175944 125424 175961
rect 140624 176175 140784 176192
rect 140624 176147 140659 176175
rect 140687 176147 140721 176175
rect 140749 176147 140784 176175
rect 140624 176113 140784 176147
rect 140624 176085 140659 176113
rect 140687 176085 140721 176113
rect 140749 176085 140784 176113
rect 140624 176051 140784 176085
rect 140624 176023 140659 176051
rect 140687 176023 140721 176051
rect 140749 176023 140784 176051
rect 140624 175989 140784 176023
rect 140624 175961 140659 175989
rect 140687 175961 140721 175989
rect 140749 175961 140784 175989
rect 140624 175944 140784 175961
rect 155984 176175 156144 176192
rect 155984 176147 156019 176175
rect 156047 176147 156081 176175
rect 156109 176147 156144 176175
rect 155984 176113 156144 176147
rect 155984 176085 156019 176113
rect 156047 176085 156081 176113
rect 156109 176085 156144 176113
rect 155984 176051 156144 176085
rect 155984 176023 156019 176051
rect 156047 176023 156081 176051
rect 156109 176023 156144 176051
rect 155984 175989 156144 176023
rect 155984 175961 156019 175989
rect 156047 175961 156081 175989
rect 156109 175961 156144 175989
rect 155984 175944 156144 175961
rect 102224 173175 102384 173192
rect 102224 173147 102259 173175
rect 102287 173147 102321 173175
rect 102349 173147 102384 173175
rect 102224 173113 102384 173147
rect 102224 173085 102259 173113
rect 102287 173085 102321 173113
rect 102349 173085 102384 173113
rect 102224 173051 102384 173085
rect 102224 173023 102259 173051
rect 102287 173023 102321 173051
rect 102349 173023 102384 173051
rect 102224 172989 102384 173023
rect 102224 172961 102259 172989
rect 102287 172961 102321 172989
rect 102349 172961 102384 172989
rect 102224 172944 102384 172961
rect 117584 173175 117744 173192
rect 117584 173147 117619 173175
rect 117647 173147 117681 173175
rect 117709 173147 117744 173175
rect 117584 173113 117744 173147
rect 117584 173085 117619 173113
rect 117647 173085 117681 173113
rect 117709 173085 117744 173113
rect 117584 173051 117744 173085
rect 117584 173023 117619 173051
rect 117647 173023 117681 173051
rect 117709 173023 117744 173051
rect 117584 172989 117744 173023
rect 117584 172961 117619 172989
rect 117647 172961 117681 172989
rect 117709 172961 117744 172989
rect 117584 172944 117744 172961
rect 132944 173175 133104 173192
rect 132944 173147 132979 173175
rect 133007 173147 133041 173175
rect 133069 173147 133104 173175
rect 132944 173113 133104 173147
rect 132944 173085 132979 173113
rect 133007 173085 133041 173113
rect 133069 173085 133104 173113
rect 132944 173051 133104 173085
rect 132944 173023 132979 173051
rect 133007 173023 133041 173051
rect 133069 173023 133104 173051
rect 132944 172989 133104 173023
rect 132944 172961 132979 172989
rect 133007 172961 133041 172989
rect 133069 172961 133104 172989
rect 132944 172944 133104 172961
rect 148304 173175 148464 173192
rect 148304 173147 148339 173175
rect 148367 173147 148401 173175
rect 148429 173147 148464 173175
rect 148304 173113 148464 173147
rect 148304 173085 148339 173113
rect 148367 173085 148401 173113
rect 148429 173085 148464 173113
rect 148304 173051 148464 173085
rect 148304 173023 148339 173051
rect 148367 173023 148401 173051
rect 148429 173023 148464 173051
rect 148304 172989 148464 173023
rect 148304 172961 148339 172989
rect 148367 172961 148401 172989
rect 148429 172961 148464 172989
rect 148304 172944 148464 172961
rect 163664 173175 163824 173192
rect 163664 173147 163699 173175
rect 163727 173147 163761 173175
rect 163789 173147 163824 173175
rect 163664 173113 163824 173147
rect 163664 173085 163699 173113
rect 163727 173085 163761 173113
rect 163789 173085 163824 173113
rect 163664 173051 163824 173085
rect 163664 173023 163699 173051
rect 163727 173023 163761 173051
rect 163789 173023 163824 173051
rect 163664 172989 163824 173023
rect 163664 172961 163699 172989
rect 163727 172961 163761 172989
rect 163789 172961 163824 172989
rect 163664 172944 163824 172961
rect 171669 173175 171979 181961
rect 171669 173147 171717 173175
rect 171745 173147 171779 173175
rect 171807 173147 171841 173175
rect 171869 173147 171903 173175
rect 171931 173147 171979 173175
rect 171669 173113 171979 173147
rect 171669 173085 171717 173113
rect 171745 173085 171779 173113
rect 171807 173085 171841 173113
rect 171869 173085 171903 173113
rect 171931 173085 171979 173113
rect 171669 173051 171979 173085
rect 171669 173023 171717 173051
rect 171745 173023 171779 173051
rect 171807 173023 171841 173051
rect 171869 173023 171903 173051
rect 171931 173023 171979 173051
rect 171669 172989 171979 173023
rect 171669 172961 171717 172989
rect 171745 172961 171779 172989
rect 171807 172961 171841 172989
rect 171869 172961 171903 172989
rect 171931 172961 171979 172989
rect 96729 167147 96777 167175
rect 96805 167147 96839 167175
rect 96867 167147 96901 167175
rect 96929 167147 96963 167175
rect 96991 167147 97039 167175
rect 96729 167113 97039 167147
rect 96729 167085 96777 167113
rect 96805 167085 96839 167113
rect 96867 167085 96901 167113
rect 96929 167085 96963 167113
rect 96991 167085 97039 167113
rect 96729 167051 97039 167085
rect 96729 167023 96777 167051
rect 96805 167023 96839 167051
rect 96867 167023 96901 167051
rect 96929 167023 96963 167051
rect 96991 167023 97039 167051
rect 96729 166989 97039 167023
rect 96729 166961 96777 166989
rect 96805 166961 96839 166989
rect 96867 166961 96901 166989
rect 96929 166961 96963 166989
rect 96991 166961 97039 166989
rect 96729 158175 97039 166961
rect 171669 164175 171979 172961
rect 171669 164147 171717 164175
rect 171745 164147 171779 164175
rect 171807 164147 171841 164175
rect 171869 164147 171903 164175
rect 171931 164147 171979 164175
rect 171669 164113 171979 164147
rect 171669 164085 171717 164113
rect 171745 164085 171779 164113
rect 171807 164085 171841 164113
rect 171869 164085 171903 164113
rect 171931 164085 171979 164113
rect 171669 164051 171979 164085
rect 171669 164023 171717 164051
rect 171745 164023 171779 164051
rect 171807 164023 171841 164051
rect 171869 164023 171903 164051
rect 171931 164023 171979 164051
rect 171669 163989 171979 164023
rect 171669 163961 171717 163989
rect 171745 163961 171779 163989
rect 171807 163961 171841 163989
rect 171869 163961 171903 163989
rect 171931 163961 171979 163989
rect 171669 158767 171979 163961
rect 173529 299086 173839 299134
rect 173529 299058 173577 299086
rect 173605 299058 173639 299086
rect 173667 299058 173701 299086
rect 173729 299058 173763 299086
rect 173791 299058 173839 299086
rect 173529 299024 173839 299058
rect 173529 298996 173577 299024
rect 173605 298996 173639 299024
rect 173667 298996 173701 299024
rect 173729 298996 173763 299024
rect 173791 298996 173839 299024
rect 173529 298962 173839 298996
rect 173529 298934 173577 298962
rect 173605 298934 173639 298962
rect 173667 298934 173701 298962
rect 173729 298934 173763 298962
rect 173791 298934 173839 298962
rect 173529 298900 173839 298934
rect 173529 298872 173577 298900
rect 173605 298872 173639 298900
rect 173667 298872 173701 298900
rect 173729 298872 173763 298900
rect 173791 298872 173839 298900
rect 173529 293175 173839 298872
rect 173529 293147 173577 293175
rect 173605 293147 173639 293175
rect 173667 293147 173701 293175
rect 173729 293147 173763 293175
rect 173791 293147 173839 293175
rect 173529 293113 173839 293147
rect 173529 293085 173577 293113
rect 173605 293085 173639 293113
rect 173667 293085 173701 293113
rect 173729 293085 173763 293113
rect 173791 293085 173839 293113
rect 173529 293051 173839 293085
rect 173529 293023 173577 293051
rect 173605 293023 173639 293051
rect 173667 293023 173701 293051
rect 173729 293023 173763 293051
rect 173791 293023 173839 293051
rect 173529 292989 173839 293023
rect 173529 292961 173577 292989
rect 173605 292961 173639 292989
rect 173667 292961 173701 292989
rect 173729 292961 173763 292989
rect 173791 292961 173839 292989
rect 173529 284175 173839 292961
rect 173529 284147 173577 284175
rect 173605 284147 173639 284175
rect 173667 284147 173701 284175
rect 173729 284147 173763 284175
rect 173791 284147 173839 284175
rect 173529 284113 173839 284147
rect 173529 284085 173577 284113
rect 173605 284085 173639 284113
rect 173667 284085 173701 284113
rect 173729 284085 173763 284113
rect 173791 284085 173839 284113
rect 173529 284051 173839 284085
rect 173529 284023 173577 284051
rect 173605 284023 173639 284051
rect 173667 284023 173701 284051
rect 173729 284023 173763 284051
rect 173791 284023 173839 284051
rect 173529 283989 173839 284023
rect 173529 283961 173577 283989
rect 173605 283961 173639 283989
rect 173667 283961 173701 283989
rect 173729 283961 173763 283989
rect 173791 283961 173839 283989
rect 173529 275175 173839 283961
rect 173529 275147 173577 275175
rect 173605 275147 173639 275175
rect 173667 275147 173701 275175
rect 173729 275147 173763 275175
rect 173791 275147 173839 275175
rect 173529 275113 173839 275147
rect 173529 275085 173577 275113
rect 173605 275085 173639 275113
rect 173667 275085 173701 275113
rect 173729 275085 173763 275113
rect 173791 275085 173839 275113
rect 173529 275051 173839 275085
rect 173529 275023 173577 275051
rect 173605 275023 173639 275051
rect 173667 275023 173701 275051
rect 173729 275023 173763 275051
rect 173791 275023 173839 275051
rect 173529 274989 173839 275023
rect 173529 274961 173577 274989
rect 173605 274961 173639 274989
rect 173667 274961 173701 274989
rect 173729 274961 173763 274989
rect 173791 274961 173839 274989
rect 173529 266175 173839 274961
rect 173529 266147 173577 266175
rect 173605 266147 173639 266175
rect 173667 266147 173701 266175
rect 173729 266147 173763 266175
rect 173791 266147 173839 266175
rect 173529 266113 173839 266147
rect 173529 266085 173577 266113
rect 173605 266085 173639 266113
rect 173667 266085 173701 266113
rect 173729 266085 173763 266113
rect 173791 266085 173839 266113
rect 173529 266051 173839 266085
rect 173529 266023 173577 266051
rect 173605 266023 173639 266051
rect 173667 266023 173701 266051
rect 173729 266023 173763 266051
rect 173791 266023 173839 266051
rect 173529 265989 173839 266023
rect 173529 265961 173577 265989
rect 173605 265961 173639 265989
rect 173667 265961 173701 265989
rect 173729 265961 173763 265989
rect 173791 265961 173839 265989
rect 173529 257175 173839 265961
rect 173529 257147 173577 257175
rect 173605 257147 173639 257175
rect 173667 257147 173701 257175
rect 173729 257147 173763 257175
rect 173791 257147 173839 257175
rect 173529 257113 173839 257147
rect 173529 257085 173577 257113
rect 173605 257085 173639 257113
rect 173667 257085 173701 257113
rect 173729 257085 173763 257113
rect 173791 257085 173839 257113
rect 173529 257051 173839 257085
rect 173529 257023 173577 257051
rect 173605 257023 173639 257051
rect 173667 257023 173701 257051
rect 173729 257023 173763 257051
rect 173791 257023 173839 257051
rect 173529 256989 173839 257023
rect 173529 256961 173577 256989
rect 173605 256961 173639 256989
rect 173667 256961 173701 256989
rect 173729 256961 173763 256989
rect 173791 256961 173839 256989
rect 173529 248175 173839 256961
rect 173529 248147 173577 248175
rect 173605 248147 173639 248175
rect 173667 248147 173701 248175
rect 173729 248147 173763 248175
rect 173791 248147 173839 248175
rect 173529 248113 173839 248147
rect 173529 248085 173577 248113
rect 173605 248085 173639 248113
rect 173667 248085 173701 248113
rect 173729 248085 173763 248113
rect 173791 248085 173839 248113
rect 173529 248051 173839 248085
rect 173529 248023 173577 248051
rect 173605 248023 173639 248051
rect 173667 248023 173701 248051
rect 173729 248023 173763 248051
rect 173791 248023 173839 248051
rect 173529 247989 173839 248023
rect 173529 247961 173577 247989
rect 173605 247961 173639 247989
rect 173667 247961 173701 247989
rect 173729 247961 173763 247989
rect 173791 247961 173839 247989
rect 173529 239175 173839 247961
rect 173529 239147 173577 239175
rect 173605 239147 173639 239175
rect 173667 239147 173701 239175
rect 173729 239147 173763 239175
rect 173791 239147 173839 239175
rect 173529 239113 173839 239147
rect 173529 239085 173577 239113
rect 173605 239085 173639 239113
rect 173667 239085 173701 239113
rect 173729 239085 173763 239113
rect 173791 239085 173839 239113
rect 173529 239051 173839 239085
rect 173529 239023 173577 239051
rect 173605 239023 173639 239051
rect 173667 239023 173701 239051
rect 173729 239023 173763 239051
rect 173791 239023 173839 239051
rect 173529 238989 173839 239023
rect 173529 238961 173577 238989
rect 173605 238961 173639 238989
rect 173667 238961 173701 238989
rect 173729 238961 173763 238989
rect 173791 238961 173839 238989
rect 173529 230175 173839 238961
rect 173529 230147 173577 230175
rect 173605 230147 173639 230175
rect 173667 230147 173701 230175
rect 173729 230147 173763 230175
rect 173791 230147 173839 230175
rect 173529 230113 173839 230147
rect 173529 230085 173577 230113
rect 173605 230085 173639 230113
rect 173667 230085 173701 230113
rect 173729 230085 173763 230113
rect 173791 230085 173839 230113
rect 173529 230051 173839 230085
rect 173529 230023 173577 230051
rect 173605 230023 173639 230051
rect 173667 230023 173701 230051
rect 173729 230023 173763 230051
rect 173791 230023 173839 230051
rect 173529 229989 173839 230023
rect 173529 229961 173577 229989
rect 173605 229961 173639 229989
rect 173667 229961 173701 229989
rect 173729 229961 173763 229989
rect 173791 229961 173839 229989
rect 173529 221175 173839 229961
rect 173529 221147 173577 221175
rect 173605 221147 173639 221175
rect 173667 221147 173701 221175
rect 173729 221147 173763 221175
rect 173791 221147 173839 221175
rect 173529 221113 173839 221147
rect 173529 221085 173577 221113
rect 173605 221085 173639 221113
rect 173667 221085 173701 221113
rect 173729 221085 173763 221113
rect 173791 221085 173839 221113
rect 173529 221051 173839 221085
rect 173529 221023 173577 221051
rect 173605 221023 173639 221051
rect 173667 221023 173701 221051
rect 173729 221023 173763 221051
rect 173791 221023 173839 221051
rect 173529 220989 173839 221023
rect 173529 220961 173577 220989
rect 173605 220961 173639 220989
rect 173667 220961 173701 220989
rect 173729 220961 173763 220989
rect 173791 220961 173839 220989
rect 173529 212175 173839 220961
rect 173529 212147 173577 212175
rect 173605 212147 173639 212175
rect 173667 212147 173701 212175
rect 173729 212147 173763 212175
rect 173791 212147 173839 212175
rect 173529 212113 173839 212147
rect 173529 212085 173577 212113
rect 173605 212085 173639 212113
rect 173667 212085 173701 212113
rect 173729 212085 173763 212113
rect 173791 212085 173839 212113
rect 173529 212051 173839 212085
rect 173529 212023 173577 212051
rect 173605 212023 173639 212051
rect 173667 212023 173701 212051
rect 173729 212023 173763 212051
rect 173791 212023 173839 212051
rect 173529 211989 173839 212023
rect 173529 211961 173577 211989
rect 173605 211961 173639 211989
rect 173667 211961 173701 211989
rect 173729 211961 173763 211989
rect 173791 211961 173839 211989
rect 173529 203175 173839 211961
rect 173529 203147 173577 203175
rect 173605 203147 173639 203175
rect 173667 203147 173701 203175
rect 173729 203147 173763 203175
rect 173791 203147 173839 203175
rect 173529 203113 173839 203147
rect 173529 203085 173577 203113
rect 173605 203085 173639 203113
rect 173667 203085 173701 203113
rect 173729 203085 173763 203113
rect 173791 203085 173839 203113
rect 173529 203051 173839 203085
rect 173529 203023 173577 203051
rect 173605 203023 173639 203051
rect 173667 203023 173701 203051
rect 173729 203023 173763 203051
rect 173791 203023 173839 203051
rect 173529 202989 173839 203023
rect 173529 202961 173577 202989
rect 173605 202961 173639 202989
rect 173667 202961 173701 202989
rect 173729 202961 173763 202989
rect 173791 202961 173839 202989
rect 173529 194175 173839 202961
rect 173529 194147 173577 194175
rect 173605 194147 173639 194175
rect 173667 194147 173701 194175
rect 173729 194147 173763 194175
rect 173791 194147 173839 194175
rect 173529 194113 173839 194147
rect 173529 194085 173577 194113
rect 173605 194085 173639 194113
rect 173667 194085 173701 194113
rect 173729 194085 173763 194113
rect 173791 194085 173839 194113
rect 173529 194051 173839 194085
rect 173529 194023 173577 194051
rect 173605 194023 173639 194051
rect 173667 194023 173701 194051
rect 173729 194023 173763 194051
rect 173791 194023 173839 194051
rect 173529 193989 173839 194023
rect 173529 193961 173577 193989
rect 173605 193961 173639 193989
rect 173667 193961 173701 193989
rect 173729 193961 173763 193989
rect 173791 193961 173839 193989
rect 173529 185175 173839 193961
rect 187029 298606 187339 299134
rect 187029 298578 187077 298606
rect 187105 298578 187139 298606
rect 187167 298578 187201 298606
rect 187229 298578 187263 298606
rect 187291 298578 187339 298606
rect 187029 298544 187339 298578
rect 187029 298516 187077 298544
rect 187105 298516 187139 298544
rect 187167 298516 187201 298544
rect 187229 298516 187263 298544
rect 187291 298516 187339 298544
rect 187029 298482 187339 298516
rect 187029 298454 187077 298482
rect 187105 298454 187139 298482
rect 187167 298454 187201 298482
rect 187229 298454 187263 298482
rect 187291 298454 187339 298482
rect 187029 298420 187339 298454
rect 187029 298392 187077 298420
rect 187105 298392 187139 298420
rect 187167 298392 187201 298420
rect 187229 298392 187263 298420
rect 187291 298392 187339 298420
rect 187029 290175 187339 298392
rect 187029 290147 187077 290175
rect 187105 290147 187139 290175
rect 187167 290147 187201 290175
rect 187229 290147 187263 290175
rect 187291 290147 187339 290175
rect 187029 290113 187339 290147
rect 187029 290085 187077 290113
rect 187105 290085 187139 290113
rect 187167 290085 187201 290113
rect 187229 290085 187263 290113
rect 187291 290085 187339 290113
rect 187029 290051 187339 290085
rect 187029 290023 187077 290051
rect 187105 290023 187139 290051
rect 187167 290023 187201 290051
rect 187229 290023 187263 290051
rect 187291 290023 187339 290051
rect 187029 289989 187339 290023
rect 187029 289961 187077 289989
rect 187105 289961 187139 289989
rect 187167 289961 187201 289989
rect 187229 289961 187263 289989
rect 187291 289961 187339 289989
rect 187029 281175 187339 289961
rect 187029 281147 187077 281175
rect 187105 281147 187139 281175
rect 187167 281147 187201 281175
rect 187229 281147 187263 281175
rect 187291 281147 187339 281175
rect 187029 281113 187339 281147
rect 187029 281085 187077 281113
rect 187105 281085 187139 281113
rect 187167 281085 187201 281113
rect 187229 281085 187263 281113
rect 187291 281085 187339 281113
rect 187029 281051 187339 281085
rect 187029 281023 187077 281051
rect 187105 281023 187139 281051
rect 187167 281023 187201 281051
rect 187229 281023 187263 281051
rect 187291 281023 187339 281051
rect 187029 280989 187339 281023
rect 187029 280961 187077 280989
rect 187105 280961 187139 280989
rect 187167 280961 187201 280989
rect 187229 280961 187263 280989
rect 187291 280961 187339 280989
rect 187029 272175 187339 280961
rect 187029 272147 187077 272175
rect 187105 272147 187139 272175
rect 187167 272147 187201 272175
rect 187229 272147 187263 272175
rect 187291 272147 187339 272175
rect 187029 272113 187339 272147
rect 187029 272085 187077 272113
rect 187105 272085 187139 272113
rect 187167 272085 187201 272113
rect 187229 272085 187263 272113
rect 187291 272085 187339 272113
rect 187029 272051 187339 272085
rect 187029 272023 187077 272051
rect 187105 272023 187139 272051
rect 187167 272023 187201 272051
rect 187229 272023 187263 272051
rect 187291 272023 187339 272051
rect 187029 271989 187339 272023
rect 187029 271961 187077 271989
rect 187105 271961 187139 271989
rect 187167 271961 187201 271989
rect 187229 271961 187263 271989
rect 187291 271961 187339 271989
rect 187029 263175 187339 271961
rect 187029 263147 187077 263175
rect 187105 263147 187139 263175
rect 187167 263147 187201 263175
rect 187229 263147 187263 263175
rect 187291 263147 187339 263175
rect 187029 263113 187339 263147
rect 187029 263085 187077 263113
rect 187105 263085 187139 263113
rect 187167 263085 187201 263113
rect 187229 263085 187263 263113
rect 187291 263085 187339 263113
rect 187029 263051 187339 263085
rect 187029 263023 187077 263051
rect 187105 263023 187139 263051
rect 187167 263023 187201 263051
rect 187229 263023 187263 263051
rect 187291 263023 187339 263051
rect 187029 262989 187339 263023
rect 187029 262961 187077 262989
rect 187105 262961 187139 262989
rect 187167 262961 187201 262989
rect 187229 262961 187263 262989
rect 187291 262961 187339 262989
rect 187029 254175 187339 262961
rect 187029 254147 187077 254175
rect 187105 254147 187139 254175
rect 187167 254147 187201 254175
rect 187229 254147 187263 254175
rect 187291 254147 187339 254175
rect 187029 254113 187339 254147
rect 187029 254085 187077 254113
rect 187105 254085 187139 254113
rect 187167 254085 187201 254113
rect 187229 254085 187263 254113
rect 187291 254085 187339 254113
rect 187029 254051 187339 254085
rect 187029 254023 187077 254051
rect 187105 254023 187139 254051
rect 187167 254023 187201 254051
rect 187229 254023 187263 254051
rect 187291 254023 187339 254051
rect 187029 253989 187339 254023
rect 187029 253961 187077 253989
rect 187105 253961 187139 253989
rect 187167 253961 187201 253989
rect 187229 253961 187263 253989
rect 187291 253961 187339 253989
rect 187029 245175 187339 253961
rect 187029 245147 187077 245175
rect 187105 245147 187139 245175
rect 187167 245147 187201 245175
rect 187229 245147 187263 245175
rect 187291 245147 187339 245175
rect 187029 245113 187339 245147
rect 187029 245085 187077 245113
rect 187105 245085 187139 245113
rect 187167 245085 187201 245113
rect 187229 245085 187263 245113
rect 187291 245085 187339 245113
rect 187029 245051 187339 245085
rect 187029 245023 187077 245051
rect 187105 245023 187139 245051
rect 187167 245023 187201 245051
rect 187229 245023 187263 245051
rect 187291 245023 187339 245051
rect 187029 244989 187339 245023
rect 187029 244961 187077 244989
rect 187105 244961 187139 244989
rect 187167 244961 187201 244989
rect 187229 244961 187263 244989
rect 187291 244961 187339 244989
rect 187029 236175 187339 244961
rect 187029 236147 187077 236175
rect 187105 236147 187139 236175
rect 187167 236147 187201 236175
rect 187229 236147 187263 236175
rect 187291 236147 187339 236175
rect 187029 236113 187339 236147
rect 187029 236085 187077 236113
rect 187105 236085 187139 236113
rect 187167 236085 187201 236113
rect 187229 236085 187263 236113
rect 187291 236085 187339 236113
rect 187029 236051 187339 236085
rect 187029 236023 187077 236051
rect 187105 236023 187139 236051
rect 187167 236023 187201 236051
rect 187229 236023 187263 236051
rect 187291 236023 187339 236051
rect 187029 235989 187339 236023
rect 187029 235961 187077 235989
rect 187105 235961 187139 235989
rect 187167 235961 187201 235989
rect 187229 235961 187263 235989
rect 187291 235961 187339 235989
rect 187029 227175 187339 235961
rect 187029 227147 187077 227175
rect 187105 227147 187139 227175
rect 187167 227147 187201 227175
rect 187229 227147 187263 227175
rect 187291 227147 187339 227175
rect 187029 227113 187339 227147
rect 187029 227085 187077 227113
rect 187105 227085 187139 227113
rect 187167 227085 187201 227113
rect 187229 227085 187263 227113
rect 187291 227085 187339 227113
rect 187029 227051 187339 227085
rect 187029 227023 187077 227051
rect 187105 227023 187139 227051
rect 187167 227023 187201 227051
rect 187229 227023 187263 227051
rect 187291 227023 187339 227051
rect 187029 226989 187339 227023
rect 187029 226961 187077 226989
rect 187105 226961 187139 226989
rect 187167 226961 187201 226989
rect 187229 226961 187263 226989
rect 187291 226961 187339 226989
rect 187029 218175 187339 226961
rect 187029 218147 187077 218175
rect 187105 218147 187139 218175
rect 187167 218147 187201 218175
rect 187229 218147 187263 218175
rect 187291 218147 187339 218175
rect 187029 218113 187339 218147
rect 187029 218085 187077 218113
rect 187105 218085 187139 218113
rect 187167 218085 187201 218113
rect 187229 218085 187263 218113
rect 187291 218085 187339 218113
rect 187029 218051 187339 218085
rect 187029 218023 187077 218051
rect 187105 218023 187139 218051
rect 187167 218023 187201 218051
rect 187229 218023 187263 218051
rect 187291 218023 187339 218051
rect 187029 217989 187339 218023
rect 187029 217961 187077 217989
rect 187105 217961 187139 217989
rect 187167 217961 187201 217989
rect 187229 217961 187263 217989
rect 187291 217961 187339 217989
rect 187029 209175 187339 217961
rect 187029 209147 187077 209175
rect 187105 209147 187139 209175
rect 187167 209147 187201 209175
rect 187229 209147 187263 209175
rect 187291 209147 187339 209175
rect 187029 209113 187339 209147
rect 187029 209085 187077 209113
rect 187105 209085 187139 209113
rect 187167 209085 187201 209113
rect 187229 209085 187263 209113
rect 187291 209085 187339 209113
rect 187029 209051 187339 209085
rect 187029 209023 187077 209051
rect 187105 209023 187139 209051
rect 187167 209023 187201 209051
rect 187229 209023 187263 209051
rect 187291 209023 187339 209051
rect 187029 208989 187339 209023
rect 187029 208961 187077 208989
rect 187105 208961 187139 208989
rect 187167 208961 187201 208989
rect 187229 208961 187263 208989
rect 187291 208961 187339 208989
rect 187029 200175 187339 208961
rect 187029 200147 187077 200175
rect 187105 200147 187139 200175
rect 187167 200147 187201 200175
rect 187229 200147 187263 200175
rect 187291 200147 187339 200175
rect 187029 200113 187339 200147
rect 187029 200085 187077 200113
rect 187105 200085 187139 200113
rect 187167 200085 187201 200113
rect 187229 200085 187263 200113
rect 187291 200085 187339 200113
rect 187029 200051 187339 200085
rect 187029 200023 187077 200051
rect 187105 200023 187139 200051
rect 187167 200023 187201 200051
rect 187229 200023 187263 200051
rect 187291 200023 187339 200051
rect 187029 199989 187339 200023
rect 187029 199961 187077 199989
rect 187105 199961 187139 199989
rect 187167 199961 187201 199989
rect 187229 199961 187263 199989
rect 187291 199961 187339 199989
rect 187029 191711 187339 199961
rect 188889 299086 189199 299134
rect 188889 299058 188937 299086
rect 188965 299058 188999 299086
rect 189027 299058 189061 299086
rect 189089 299058 189123 299086
rect 189151 299058 189199 299086
rect 188889 299024 189199 299058
rect 188889 298996 188937 299024
rect 188965 298996 188999 299024
rect 189027 298996 189061 299024
rect 189089 298996 189123 299024
rect 189151 298996 189199 299024
rect 188889 298962 189199 298996
rect 188889 298934 188937 298962
rect 188965 298934 188999 298962
rect 189027 298934 189061 298962
rect 189089 298934 189123 298962
rect 189151 298934 189199 298962
rect 188889 298900 189199 298934
rect 188889 298872 188937 298900
rect 188965 298872 188999 298900
rect 189027 298872 189061 298900
rect 189089 298872 189123 298900
rect 189151 298872 189199 298900
rect 188889 293175 189199 298872
rect 188889 293147 188937 293175
rect 188965 293147 188999 293175
rect 189027 293147 189061 293175
rect 189089 293147 189123 293175
rect 189151 293147 189199 293175
rect 188889 293113 189199 293147
rect 188889 293085 188937 293113
rect 188965 293085 188999 293113
rect 189027 293085 189061 293113
rect 189089 293085 189123 293113
rect 189151 293085 189199 293113
rect 188889 293051 189199 293085
rect 188889 293023 188937 293051
rect 188965 293023 188999 293051
rect 189027 293023 189061 293051
rect 189089 293023 189123 293051
rect 189151 293023 189199 293051
rect 188889 292989 189199 293023
rect 188889 292961 188937 292989
rect 188965 292961 188999 292989
rect 189027 292961 189061 292989
rect 189089 292961 189123 292989
rect 189151 292961 189199 292989
rect 188889 284175 189199 292961
rect 188889 284147 188937 284175
rect 188965 284147 188999 284175
rect 189027 284147 189061 284175
rect 189089 284147 189123 284175
rect 189151 284147 189199 284175
rect 188889 284113 189199 284147
rect 188889 284085 188937 284113
rect 188965 284085 188999 284113
rect 189027 284085 189061 284113
rect 189089 284085 189123 284113
rect 189151 284085 189199 284113
rect 188889 284051 189199 284085
rect 188889 284023 188937 284051
rect 188965 284023 188999 284051
rect 189027 284023 189061 284051
rect 189089 284023 189123 284051
rect 189151 284023 189199 284051
rect 188889 283989 189199 284023
rect 188889 283961 188937 283989
rect 188965 283961 188999 283989
rect 189027 283961 189061 283989
rect 189089 283961 189123 283989
rect 189151 283961 189199 283989
rect 188889 275175 189199 283961
rect 188889 275147 188937 275175
rect 188965 275147 188999 275175
rect 189027 275147 189061 275175
rect 189089 275147 189123 275175
rect 189151 275147 189199 275175
rect 188889 275113 189199 275147
rect 188889 275085 188937 275113
rect 188965 275085 188999 275113
rect 189027 275085 189061 275113
rect 189089 275085 189123 275113
rect 189151 275085 189199 275113
rect 188889 275051 189199 275085
rect 188889 275023 188937 275051
rect 188965 275023 188999 275051
rect 189027 275023 189061 275051
rect 189089 275023 189123 275051
rect 189151 275023 189199 275051
rect 188889 274989 189199 275023
rect 188889 274961 188937 274989
rect 188965 274961 188999 274989
rect 189027 274961 189061 274989
rect 189089 274961 189123 274989
rect 189151 274961 189199 274989
rect 188889 266175 189199 274961
rect 188889 266147 188937 266175
rect 188965 266147 188999 266175
rect 189027 266147 189061 266175
rect 189089 266147 189123 266175
rect 189151 266147 189199 266175
rect 188889 266113 189199 266147
rect 188889 266085 188937 266113
rect 188965 266085 188999 266113
rect 189027 266085 189061 266113
rect 189089 266085 189123 266113
rect 189151 266085 189199 266113
rect 188889 266051 189199 266085
rect 188889 266023 188937 266051
rect 188965 266023 188999 266051
rect 189027 266023 189061 266051
rect 189089 266023 189123 266051
rect 189151 266023 189199 266051
rect 188889 265989 189199 266023
rect 188889 265961 188937 265989
rect 188965 265961 188999 265989
rect 189027 265961 189061 265989
rect 189089 265961 189123 265989
rect 189151 265961 189199 265989
rect 188889 257175 189199 265961
rect 188889 257147 188937 257175
rect 188965 257147 188999 257175
rect 189027 257147 189061 257175
rect 189089 257147 189123 257175
rect 189151 257147 189199 257175
rect 188889 257113 189199 257147
rect 188889 257085 188937 257113
rect 188965 257085 188999 257113
rect 189027 257085 189061 257113
rect 189089 257085 189123 257113
rect 189151 257085 189199 257113
rect 188889 257051 189199 257085
rect 188889 257023 188937 257051
rect 188965 257023 188999 257051
rect 189027 257023 189061 257051
rect 189089 257023 189123 257051
rect 189151 257023 189199 257051
rect 188889 256989 189199 257023
rect 188889 256961 188937 256989
rect 188965 256961 188999 256989
rect 189027 256961 189061 256989
rect 189089 256961 189123 256989
rect 189151 256961 189199 256989
rect 188889 248175 189199 256961
rect 188889 248147 188937 248175
rect 188965 248147 188999 248175
rect 189027 248147 189061 248175
rect 189089 248147 189123 248175
rect 189151 248147 189199 248175
rect 188889 248113 189199 248147
rect 188889 248085 188937 248113
rect 188965 248085 188999 248113
rect 189027 248085 189061 248113
rect 189089 248085 189123 248113
rect 189151 248085 189199 248113
rect 188889 248051 189199 248085
rect 188889 248023 188937 248051
rect 188965 248023 188999 248051
rect 189027 248023 189061 248051
rect 189089 248023 189123 248051
rect 189151 248023 189199 248051
rect 188889 247989 189199 248023
rect 188889 247961 188937 247989
rect 188965 247961 188999 247989
rect 189027 247961 189061 247989
rect 189089 247961 189123 247989
rect 189151 247961 189199 247989
rect 188889 239175 189199 247961
rect 188889 239147 188937 239175
rect 188965 239147 188999 239175
rect 189027 239147 189061 239175
rect 189089 239147 189123 239175
rect 189151 239147 189199 239175
rect 188889 239113 189199 239147
rect 188889 239085 188937 239113
rect 188965 239085 188999 239113
rect 189027 239085 189061 239113
rect 189089 239085 189123 239113
rect 189151 239085 189199 239113
rect 188889 239051 189199 239085
rect 188889 239023 188937 239051
rect 188965 239023 188999 239051
rect 189027 239023 189061 239051
rect 189089 239023 189123 239051
rect 189151 239023 189199 239051
rect 188889 238989 189199 239023
rect 188889 238961 188937 238989
rect 188965 238961 188999 238989
rect 189027 238961 189061 238989
rect 189089 238961 189123 238989
rect 189151 238961 189199 238989
rect 188889 230175 189199 238961
rect 188889 230147 188937 230175
rect 188965 230147 188999 230175
rect 189027 230147 189061 230175
rect 189089 230147 189123 230175
rect 189151 230147 189199 230175
rect 188889 230113 189199 230147
rect 188889 230085 188937 230113
rect 188965 230085 188999 230113
rect 189027 230085 189061 230113
rect 189089 230085 189123 230113
rect 189151 230085 189199 230113
rect 188889 230051 189199 230085
rect 188889 230023 188937 230051
rect 188965 230023 188999 230051
rect 189027 230023 189061 230051
rect 189089 230023 189123 230051
rect 189151 230023 189199 230051
rect 188889 229989 189199 230023
rect 188889 229961 188937 229989
rect 188965 229961 188999 229989
rect 189027 229961 189061 229989
rect 189089 229961 189123 229989
rect 189151 229961 189199 229989
rect 188889 221175 189199 229961
rect 188889 221147 188937 221175
rect 188965 221147 188999 221175
rect 189027 221147 189061 221175
rect 189089 221147 189123 221175
rect 189151 221147 189199 221175
rect 188889 221113 189199 221147
rect 188889 221085 188937 221113
rect 188965 221085 188999 221113
rect 189027 221085 189061 221113
rect 189089 221085 189123 221113
rect 189151 221085 189199 221113
rect 188889 221051 189199 221085
rect 188889 221023 188937 221051
rect 188965 221023 188999 221051
rect 189027 221023 189061 221051
rect 189089 221023 189123 221051
rect 189151 221023 189199 221051
rect 188889 220989 189199 221023
rect 188889 220961 188937 220989
rect 188965 220961 188999 220989
rect 189027 220961 189061 220989
rect 189089 220961 189123 220989
rect 189151 220961 189199 220989
rect 188889 212175 189199 220961
rect 188889 212147 188937 212175
rect 188965 212147 188999 212175
rect 189027 212147 189061 212175
rect 189089 212147 189123 212175
rect 189151 212147 189199 212175
rect 188889 212113 189199 212147
rect 188889 212085 188937 212113
rect 188965 212085 188999 212113
rect 189027 212085 189061 212113
rect 189089 212085 189123 212113
rect 189151 212085 189199 212113
rect 188889 212051 189199 212085
rect 188889 212023 188937 212051
rect 188965 212023 188999 212051
rect 189027 212023 189061 212051
rect 189089 212023 189123 212051
rect 189151 212023 189199 212051
rect 188889 211989 189199 212023
rect 188889 211961 188937 211989
rect 188965 211961 188999 211989
rect 189027 211961 189061 211989
rect 189089 211961 189123 211989
rect 189151 211961 189199 211989
rect 188889 203175 189199 211961
rect 188889 203147 188937 203175
rect 188965 203147 188999 203175
rect 189027 203147 189061 203175
rect 189089 203147 189123 203175
rect 189151 203147 189199 203175
rect 188889 203113 189199 203147
rect 188889 203085 188937 203113
rect 188965 203085 188999 203113
rect 189027 203085 189061 203113
rect 189089 203085 189123 203113
rect 189151 203085 189199 203113
rect 188889 203051 189199 203085
rect 188889 203023 188937 203051
rect 188965 203023 188999 203051
rect 189027 203023 189061 203051
rect 189089 203023 189123 203051
rect 189151 203023 189199 203051
rect 188889 202989 189199 203023
rect 188889 202961 188937 202989
rect 188965 202961 188999 202989
rect 189027 202961 189061 202989
rect 189089 202961 189123 202989
rect 189151 202961 189199 202989
rect 188889 194175 189199 202961
rect 202389 298606 202699 299134
rect 202389 298578 202437 298606
rect 202465 298578 202499 298606
rect 202527 298578 202561 298606
rect 202589 298578 202623 298606
rect 202651 298578 202699 298606
rect 202389 298544 202699 298578
rect 202389 298516 202437 298544
rect 202465 298516 202499 298544
rect 202527 298516 202561 298544
rect 202589 298516 202623 298544
rect 202651 298516 202699 298544
rect 202389 298482 202699 298516
rect 202389 298454 202437 298482
rect 202465 298454 202499 298482
rect 202527 298454 202561 298482
rect 202589 298454 202623 298482
rect 202651 298454 202699 298482
rect 202389 298420 202699 298454
rect 202389 298392 202437 298420
rect 202465 298392 202499 298420
rect 202527 298392 202561 298420
rect 202589 298392 202623 298420
rect 202651 298392 202699 298420
rect 202389 290175 202699 298392
rect 202389 290147 202437 290175
rect 202465 290147 202499 290175
rect 202527 290147 202561 290175
rect 202589 290147 202623 290175
rect 202651 290147 202699 290175
rect 202389 290113 202699 290147
rect 202389 290085 202437 290113
rect 202465 290085 202499 290113
rect 202527 290085 202561 290113
rect 202589 290085 202623 290113
rect 202651 290085 202699 290113
rect 202389 290051 202699 290085
rect 202389 290023 202437 290051
rect 202465 290023 202499 290051
rect 202527 290023 202561 290051
rect 202589 290023 202623 290051
rect 202651 290023 202699 290051
rect 202389 289989 202699 290023
rect 202389 289961 202437 289989
rect 202465 289961 202499 289989
rect 202527 289961 202561 289989
rect 202589 289961 202623 289989
rect 202651 289961 202699 289989
rect 202389 281175 202699 289961
rect 202389 281147 202437 281175
rect 202465 281147 202499 281175
rect 202527 281147 202561 281175
rect 202589 281147 202623 281175
rect 202651 281147 202699 281175
rect 202389 281113 202699 281147
rect 202389 281085 202437 281113
rect 202465 281085 202499 281113
rect 202527 281085 202561 281113
rect 202589 281085 202623 281113
rect 202651 281085 202699 281113
rect 202389 281051 202699 281085
rect 202389 281023 202437 281051
rect 202465 281023 202499 281051
rect 202527 281023 202561 281051
rect 202589 281023 202623 281051
rect 202651 281023 202699 281051
rect 202389 280989 202699 281023
rect 202389 280961 202437 280989
rect 202465 280961 202499 280989
rect 202527 280961 202561 280989
rect 202589 280961 202623 280989
rect 202651 280961 202699 280989
rect 202389 272175 202699 280961
rect 202389 272147 202437 272175
rect 202465 272147 202499 272175
rect 202527 272147 202561 272175
rect 202589 272147 202623 272175
rect 202651 272147 202699 272175
rect 202389 272113 202699 272147
rect 202389 272085 202437 272113
rect 202465 272085 202499 272113
rect 202527 272085 202561 272113
rect 202589 272085 202623 272113
rect 202651 272085 202699 272113
rect 202389 272051 202699 272085
rect 202389 272023 202437 272051
rect 202465 272023 202499 272051
rect 202527 272023 202561 272051
rect 202589 272023 202623 272051
rect 202651 272023 202699 272051
rect 202389 271989 202699 272023
rect 202389 271961 202437 271989
rect 202465 271961 202499 271989
rect 202527 271961 202561 271989
rect 202589 271961 202623 271989
rect 202651 271961 202699 271989
rect 202389 263175 202699 271961
rect 202389 263147 202437 263175
rect 202465 263147 202499 263175
rect 202527 263147 202561 263175
rect 202589 263147 202623 263175
rect 202651 263147 202699 263175
rect 202389 263113 202699 263147
rect 202389 263085 202437 263113
rect 202465 263085 202499 263113
rect 202527 263085 202561 263113
rect 202589 263085 202623 263113
rect 202651 263085 202699 263113
rect 202389 263051 202699 263085
rect 202389 263023 202437 263051
rect 202465 263023 202499 263051
rect 202527 263023 202561 263051
rect 202589 263023 202623 263051
rect 202651 263023 202699 263051
rect 202389 262989 202699 263023
rect 202389 262961 202437 262989
rect 202465 262961 202499 262989
rect 202527 262961 202561 262989
rect 202589 262961 202623 262989
rect 202651 262961 202699 262989
rect 202389 254175 202699 262961
rect 202389 254147 202437 254175
rect 202465 254147 202499 254175
rect 202527 254147 202561 254175
rect 202589 254147 202623 254175
rect 202651 254147 202699 254175
rect 202389 254113 202699 254147
rect 202389 254085 202437 254113
rect 202465 254085 202499 254113
rect 202527 254085 202561 254113
rect 202589 254085 202623 254113
rect 202651 254085 202699 254113
rect 202389 254051 202699 254085
rect 202389 254023 202437 254051
rect 202465 254023 202499 254051
rect 202527 254023 202561 254051
rect 202589 254023 202623 254051
rect 202651 254023 202699 254051
rect 202389 253989 202699 254023
rect 202389 253961 202437 253989
rect 202465 253961 202499 253989
rect 202527 253961 202561 253989
rect 202589 253961 202623 253989
rect 202651 253961 202699 253989
rect 202389 245175 202699 253961
rect 202389 245147 202437 245175
rect 202465 245147 202499 245175
rect 202527 245147 202561 245175
rect 202589 245147 202623 245175
rect 202651 245147 202699 245175
rect 202389 245113 202699 245147
rect 202389 245085 202437 245113
rect 202465 245085 202499 245113
rect 202527 245085 202561 245113
rect 202589 245085 202623 245113
rect 202651 245085 202699 245113
rect 202389 245051 202699 245085
rect 202389 245023 202437 245051
rect 202465 245023 202499 245051
rect 202527 245023 202561 245051
rect 202589 245023 202623 245051
rect 202651 245023 202699 245051
rect 202389 244989 202699 245023
rect 202389 244961 202437 244989
rect 202465 244961 202499 244989
rect 202527 244961 202561 244989
rect 202589 244961 202623 244989
rect 202651 244961 202699 244989
rect 202389 236175 202699 244961
rect 202389 236147 202437 236175
rect 202465 236147 202499 236175
rect 202527 236147 202561 236175
rect 202589 236147 202623 236175
rect 202651 236147 202699 236175
rect 202389 236113 202699 236147
rect 202389 236085 202437 236113
rect 202465 236085 202499 236113
rect 202527 236085 202561 236113
rect 202589 236085 202623 236113
rect 202651 236085 202699 236113
rect 202389 236051 202699 236085
rect 202389 236023 202437 236051
rect 202465 236023 202499 236051
rect 202527 236023 202561 236051
rect 202589 236023 202623 236051
rect 202651 236023 202699 236051
rect 202389 235989 202699 236023
rect 202389 235961 202437 235989
rect 202465 235961 202499 235989
rect 202527 235961 202561 235989
rect 202589 235961 202623 235989
rect 202651 235961 202699 235989
rect 202389 227175 202699 235961
rect 202389 227147 202437 227175
rect 202465 227147 202499 227175
rect 202527 227147 202561 227175
rect 202589 227147 202623 227175
rect 202651 227147 202699 227175
rect 202389 227113 202699 227147
rect 202389 227085 202437 227113
rect 202465 227085 202499 227113
rect 202527 227085 202561 227113
rect 202589 227085 202623 227113
rect 202651 227085 202699 227113
rect 202389 227051 202699 227085
rect 202389 227023 202437 227051
rect 202465 227023 202499 227051
rect 202527 227023 202561 227051
rect 202589 227023 202623 227051
rect 202651 227023 202699 227051
rect 202389 226989 202699 227023
rect 202389 226961 202437 226989
rect 202465 226961 202499 226989
rect 202527 226961 202561 226989
rect 202589 226961 202623 226989
rect 202651 226961 202699 226989
rect 202389 218175 202699 226961
rect 202389 218147 202437 218175
rect 202465 218147 202499 218175
rect 202527 218147 202561 218175
rect 202589 218147 202623 218175
rect 202651 218147 202699 218175
rect 202389 218113 202699 218147
rect 202389 218085 202437 218113
rect 202465 218085 202499 218113
rect 202527 218085 202561 218113
rect 202589 218085 202623 218113
rect 202651 218085 202699 218113
rect 202389 218051 202699 218085
rect 202389 218023 202437 218051
rect 202465 218023 202499 218051
rect 202527 218023 202561 218051
rect 202589 218023 202623 218051
rect 202651 218023 202699 218051
rect 202389 217989 202699 218023
rect 202389 217961 202437 217989
rect 202465 217961 202499 217989
rect 202527 217961 202561 217989
rect 202589 217961 202623 217989
rect 202651 217961 202699 217989
rect 202389 209175 202699 217961
rect 202389 209147 202437 209175
rect 202465 209147 202499 209175
rect 202527 209147 202561 209175
rect 202589 209147 202623 209175
rect 202651 209147 202699 209175
rect 202389 209113 202699 209147
rect 202389 209085 202437 209113
rect 202465 209085 202499 209113
rect 202527 209085 202561 209113
rect 202589 209085 202623 209113
rect 202651 209085 202699 209113
rect 202389 209051 202699 209085
rect 202389 209023 202437 209051
rect 202465 209023 202499 209051
rect 202527 209023 202561 209051
rect 202589 209023 202623 209051
rect 202651 209023 202699 209051
rect 202389 208989 202699 209023
rect 202389 208961 202437 208989
rect 202465 208961 202499 208989
rect 202527 208961 202561 208989
rect 202589 208961 202623 208989
rect 202651 208961 202699 208989
rect 202389 200175 202699 208961
rect 202389 200147 202437 200175
rect 202465 200147 202499 200175
rect 202527 200147 202561 200175
rect 202589 200147 202623 200175
rect 202651 200147 202699 200175
rect 202389 200113 202699 200147
rect 202389 200085 202437 200113
rect 202465 200085 202499 200113
rect 202527 200085 202561 200113
rect 202589 200085 202623 200113
rect 202651 200085 202699 200113
rect 202389 200051 202699 200085
rect 202389 200023 202437 200051
rect 202465 200023 202499 200051
rect 202527 200023 202561 200051
rect 202589 200023 202623 200051
rect 202651 200023 202699 200051
rect 202389 199989 202699 200023
rect 202389 199961 202437 199989
rect 202465 199961 202499 199989
rect 202527 199961 202561 199989
rect 202589 199961 202623 199989
rect 202651 199961 202699 199989
rect 188889 194147 188937 194175
rect 188965 194147 188999 194175
rect 189027 194147 189061 194175
rect 189089 194147 189123 194175
rect 189151 194147 189199 194175
rect 188889 194113 189199 194147
rect 188889 194085 188937 194113
rect 188965 194085 188999 194113
rect 189027 194085 189061 194113
rect 189089 194085 189123 194113
rect 189151 194085 189199 194113
rect 188889 194051 189199 194085
rect 188889 194023 188937 194051
rect 188965 194023 188999 194051
rect 189027 194023 189061 194051
rect 189089 194023 189123 194051
rect 189151 194023 189199 194051
rect 188889 193989 189199 194023
rect 188889 193961 188937 193989
rect 188965 193961 188999 193989
rect 189027 193961 189061 193989
rect 189089 193961 189123 193989
rect 189151 193961 189199 193989
rect 188889 191711 189199 193961
rect 189904 194175 190064 194192
rect 189904 194147 189939 194175
rect 189967 194147 190001 194175
rect 190029 194147 190064 194175
rect 189904 194113 190064 194147
rect 189904 194085 189939 194113
rect 189967 194085 190001 194113
rect 190029 194085 190064 194113
rect 189904 194051 190064 194085
rect 189904 194023 189939 194051
rect 189967 194023 190001 194051
rect 190029 194023 190064 194051
rect 189904 193989 190064 194023
rect 189904 193961 189939 193989
rect 189967 193961 190001 193989
rect 190029 193961 190064 193989
rect 189904 193944 190064 193961
rect 182224 191175 182384 191192
rect 182224 191147 182259 191175
rect 182287 191147 182321 191175
rect 182349 191147 182384 191175
rect 182224 191113 182384 191147
rect 182224 191085 182259 191113
rect 182287 191085 182321 191113
rect 182349 191085 182384 191113
rect 182224 191051 182384 191085
rect 182224 191023 182259 191051
rect 182287 191023 182321 191051
rect 182349 191023 182384 191051
rect 182224 190989 182384 191023
rect 182224 190961 182259 190989
rect 182287 190961 182321 190989
rect 182349 190961 182384 190989
rect 182224 190944 182384 190961
rect 197584 191175 197744 191192
rect 197584 191147 197619 191175
rect 197647 191147 197681 191175
rect 197709 191147 197744 191175
rect 197584 191113 197744 191147
rect 197584 191085 197619 191113
rect 197647 191085 197681 191113
rect 197709 191085 197744 191113
rect 197584 191051 197744 191085
rect 197584 191023 197619 191051
rect 197647 191023 197681 191051
rect 197709 191023 197744 191051
rect 197584 190989 197744 191023
rect 197584 190961 197619 190989
rect 197647 190961 197681 190989
rect 197709 190961 197744 190989
rect 197584 190944 197744 190961
rect 202389 191175 202699 199961
rect 202389 191147 202437 191175
rect 202465 191147 202499 191175
rect 202527 191147 202561 191175
rect 202589 191147 202623 191175
rect 202651 191147 202699 191175
rect 202389 191113 202699 191147
rect 202389 191085 202437 191113
rect 202465 191085 202499 191113
rect 202527 191085 202561 191113
rect 202589 191085 202623 191113
rect 202651 191085 202699 191113
rect 202389 191051 202699 191085
rect 202389 191023 202437 191051
rect 202465 191023 202499 191051
rect 202527 191023 202561 191051
rect 202589 191023 202623 191051
rect 202651 191023 202699 191051
rect 202389 190989 202699 191023
rect 202389 190961 202437 190989
rect 202465 190961 202499 190989
rect 202527 190961 202561 190989
rect 202589 190961 202623 190989
rect 202651 190961 202699 190989
rect 173529 185147 173577 185175
rect 173605 185147 173639 185175
rect 173667 185147 173701 185175
rect 173729 185147 173763 185175
rect 173791 185147 173839 185175
rect 173529 185113 173839 185147
rect 173529 185085 173577 185113
rect 173605 185085 173639 185113
rect 173667 185085 173701 185113
rect 173729 185085 173763 185113
rect 173791 185085 173839 185113
rect 173529 185051 173839 185085
rect 173529 185023 173577 185051
rect 173605 185023 173639 185051
rect 173667 185023 173701 185051
rect 173729 185023 173763 185051
rect 173791 185023 173839 185051
rect 173529 184989 173839 185023
rect 173529 184961 173577 184989
rect 173605 184961 173639 184989
rect 173667 184961 173701 184989
rect 173729 184961 173763 184989
rect 173791 184961 173839 184989
rect 173529 176175 173839 184961
rect 189904 185175 190064 185192
rect 189904 185147 189939 185175
rect 189967 185147 190001 185175
rect 190029 185147 190064 185175
rect 189904 185113 190064 185147
rect 189904 185085 189939 185113
rect 189967 185085 190001 185113
rect 190029 185085 190064 185113
rect 189904 185051 190064 185085
rect 189904 185023 189939 185051
rect 189967 185023 190001 185051
rect 190029 185023 190064 185051
rect 189904 184989 190064 185023
rect 189904 184961 189939 184989
rect 189967 184961 190001 184989
rect 190029 184961 190064 184989
rect 189904 184944 190064 184961
rect 182224 182175 182384 182192
rect 182224 182147 182259 182175
rect 182287 182147 182321 182175
rect 182349 182147 182384 182175
rect 182224 182113 182384 182147
rect 182224 182085 182259 182113
rect 182287 182085 182321 182113
rect 182349 182085 182384 182113
rect 182224 182051 182384 182085
rect 182224 182023 182259 182051
rect 182287 182023 182321 182051
rect 182349 182023 182384 182051
rect 182224 181989 182384 182023
rect 182224 181961 182259 181989
rect 182287 181961 182321 181989
rect 182349 181961 182384 181989
rect 182224 181944 182384 181961
rect 197584 182175 197744 182192
rect 197584 182147 197619 182175
rect 197647 182147 197681 182175
rect 197709 182147 197744 182175
rect 197584 182113 197744 182147
rect 197584 182085 197619 182113
rect 197647 182085 197681 182113
rect 197709 182085 197744 182113
rect 197584 182051 197744 182085
rect 197584 182023 197619 182051
rect 197647 182023 197681 182051
rect 197709 182023 197744 182051
rect 197584 181989 197744 182023
rect 197584 181961 197619 181989
rect 197647 181961 197681 181989
rect 197709 181961 197744 181989
rect 197584 181944 197744 181961
rect 202389 182175 202699 190961
rect 202389 182147 202437 182175
rect 202465 182147 202499 182175
rect 202527 182147 202561 182175
rect 202589 182147 202623 182175
rect 202651 182147 202699 182175
rect 202389 182113 202699 182147
rect 202389 182085 202437 182113
rect 202465 182085 202499 182113
rect 202527 182085 202561 182113
rect 202589 182085 202623 182113
rect 202651 182085 202699 182113
rect 202389 182051 202699 182085
rect 202389 182023 202437 182051
rect 202465 182023 202499 182051
rect 202527 182023 202561 182051
rect 202589 182023 202623 182051
rect 202651 182023 202699 182051
rect 202389 181989 202699 182023
rect 202389 181961 202437 181989
rect 202465 181961 202499 181989
rect 202527 181961 202561 181989
rect 202589 181961 202623 181989
rect 202651 181961 202699 181989
rect 173529 176147 173577 176175
rect 173605 176147 173639 176175
rect 173667 176147 173701 176175
rect 173729 176147 173763 176175
rect 173791 176147 173839 176175
rect 173529 176113 173839 176147
rect 173529 176085 173577 176113
rect 173605 176085 173639 176113
rect 173667 176085 173701 176113
rect 173729 176085 173763 176113
rect 173791 176085 173839 176113
rect 173529 176051 173839 176085
rect 173529 176023 173577 176051
rect 173605 176023 173639 176051
rect 173667 176023 173701 176051
rect 173729 176023 173763 176051
rect 173791 176023 173839 176051
rect 173529 175989 173839 176023
rect 173529 175961 173577 175989
rect 173605 175961 173639 175989
rect 173667 175961 173701 175989
rect 173729 175961 173763 175989
rect 173791 175961 173839 175989
rect 173529 167175 173839 175961
rect 189904 176175 190064 176192
rect 189904 176147 189939 176175
rect 189967 176147 190001 176175
rect 190029 176147 190064 176175
rect 189904 176113 190064 176147
rect 189904 176085 189939 176113
rect 189967 176085 190001 176113
rect 190029 176085 190064 176113
rect 189904 176051 190064 176085
rect 189904 176023 189939 176051
rect 189967 176023 190001 176051
rect 190029 176023 190064 176051
rect 189904 175989 190064 176023
rect 189904 175961 189939 175989
rect 189967 175961 190001 175989
rect 190029 175961 190064 175989
rect 189904 175944 190064 175961
rect 182224 173175 182384 173192
rect 182224 173147 182259 173175
rect 182287 173147 182321 173175
rect 182349 173147 182384 173175
rect 182224 173113 182384 173147
rect 182224 173085 182259 173113
rect 182287 173085 182321 173113
rect 182349 173085 182384 173113
rect 182224 173051 182384 173085
rect 182224 173023 182259 173051
rect 182287 173023 182321 173051
rect 182349 173023 182384 173051
rect 182224 172989 182384 173023
rect 182224 172961 182259 172989
rect 182287 172961 182321 172989
rect 182349 172961 182384 172989
rect 182224 172944 182384 172961
rect 187029 173175 187339 174889
rect 187029 173147 187077 173175
rect 187105 173147 187139 173175
rect 187167 173147 187201 173175
rect 187229 173147 187263 173175
rect 187291 173147 187339 173175
rect 187029 173113 187339 173147
rect 187029 173085 187077 173113
rect 187105 173085 187139 173113
rect 187167 173085 187201 173113
rect 187229 173085 187263 173113
rect 187291 173085 187339 173113
rect 187029 173051 187339 173085
rect 187029 173023 187077 173051
rect 187105 173023 187139 173051
rect 187167 173023 187201 173051
rect 187229 173023 187263 173051
rect 187291 173023 187339 173051
rect 187029 172989 187339 173023
rect 187029 172961 187077 172989
rect 187105 172961 187139 172989
rect 187167 172961 187201 172989
rect 187229 172961 187263 172989
rect 187291 172961 187339 172989
rect 173529 167147 173577 167175
rect 173605 167147 173639 167175
rect 173667 167147 173701 167175
rect 173729 167147 173763 167175
rect 173791 167147 173839 167175
rect 173529 167113 173839 167147
rect 173529 167085 173577 167113
rect 173605 167085 173639 167113
rect 173667 167085 173701 167113
rect 173729 167085 173763 167113
rect 173791 167085 173839 167113
rect 173529 167051 173839 167085
rect 173529 167023 173577 167051
rect 173605 167023 173639 167051
rect 173667 167023 173701 167051
rect 173729 167023 173763 167051
rect 173791 167023 173839 167051
rect 173529 166989 173839 167023
rect 173529 166961 173577 166989
rect 173605 166961 173639 166989
rect 173667 166961 173701 166989
rect 173729 166961 173763 166989
rect 173791 166961 173839 166989
rect 173529 158767 173839 166961
rect 187029 164175 187339 172961
rect 197584 173175 197744 173192
rect 197584 173147 197619 173175
rect 197647 173147 197681 173175
rect 197709 173147 197744 173175
rect 197584 173113 197744 173147
rect 197584 173085 197619 173113
rect 197647 173085 197681 173113
rect 197709 173085 197744 173113
rect 197584 173051 197744 173085
rect 197584 173023 197619 173051
rect 197647 173023 197681 173051
rect 197709 173023 197744 173051
rect 197584 172989 197744 173023
rect 197584 172961 197619 172989
rect 197647 172961 197681 172989
rect 197709 172961 197744 172989
rect 197584 172944 197744 172961
rect 202389 173175 202699 181961
rect 202389 173147 202437 173175
rect 202465 173147 202499 173175
rect 202527 173147 202561 173175
rect 202589 173147 202623 173175
rect 202651 173147 202699 173175
rect 202389 173113 202699 173147
rect 202389 173085 202437 173113
rect 202465 173085 202499 173113
rect 202527 173085 202561 173113
rect 202589 173085 202623 173113
rect 202651 173085 202699 173113
rect 202389 173051 202699 173085
rect 202389 173023 202437 173051
rect 202465 173023 202499 173051
rect 202527 173023 202561 173051
rect 202589 173023 202623 173051
rect 202651 173023 202699 173051
rect 202389 172989 202699 173023
rect 202389 172961 202437 172989
rect 202465 172961 202499 172989
rect 202527 172961 202561 172989
rect 202589 172961 202623 172989
rect 202651 172961 202699 172989
rect 187029 164147 187077 164175
rect 187105 164147 187139 164175
rect 187167 164147 187201 164175
rect 187229 164147 187263 164175
rect 187291 164147 187339 164175
rect 187029 164113 187339 164147
rect 187029 164085 187077 164113
rect 187105 164085 187139 164113
rect 187167 164085 187201 164113
rect 187229 164085 187263 164113
rect 187291 164085 187339 164113
rect 187029 164051 187339 164085
rect 187029 164023 187077 164051
rect 187105 164023 187139 164051
rect 187167 164023 187201 164051
rect 187229 164023 187263 164051
rect 187291 164023 187339 164051
rect 187029 163989 187339 164023
rect 187029 163961 187077 163989
rect 187105 163961 187139 163989
rect 187167 163961 187201 163989
rect 187229 163961 187263 163989
rect 187291 163961 187339 163989
rect 187029 158767 187339 163961
rect 202389 164175 202699 172961
rect 202389 164147 202437 164175
rect 202465 164147 202499 164175
rect 202527 164147 202561 164175
rect 202589 164147 202623 164175
rect 202651 164147 202699 164175
rect 202389 164113 202699 164147
rect 202389 164085 202437 164113
rect 202465 164085 202499 164113
rect 202527 164085 202561 164113
rect 202589 164085 202623 164113
rect 202651 164085 202699 164113
rect 202389 164051 202699 164085
rect 202389 164023 202437 164051
rect 202465 164023 202499 164051
rect 202527 164023 202561 164051
rect 202589 164023 202623 164051
rect 202651 164023 202699 164051
rect 202389 163989 202699 164023
rect 202389 163961 202437 163989
rect 202465 163961 202499 163989
rect 202527 163961 202561 163989
rect 202589 163961 202623 163989
rect 202651 163961 202699 163989
rect 202389 158767 202699 163961
rect 204249 299086 204559 299134
rect 204249 299058 204297 299086
rect 204325 299058 204359 299086
rect 204387 299058 204421 299086
rect 204449 299058 204483 299086
rect 204511 299058 204559 299086
rect 204249 299024 204559 299058
rect 204249 298996 204297 299024
rect 204325 298996 204359 299024
rect 204387 298996 204421 299024
rect 204449 298996 204483 299024
rect 204511 298996 204559 299024
rect 204249 298962 204559 298996
rect 204249 298934 204297 298962
rect 204325 298934 204359 298962
rect 204387 298934 204421 298962
rect 204449 298934 204483 298962
rect 204511 298934 204559 298962
rect 204249 298900 204559 298934
rect 204249 298872 204297 298900
rect 204325 298872 204359 298900
rect 204387 298872 204421 298900
rect 204449 298872 204483 298900
rect 204511 298872 204559 298900
rect 204249 293175 204559 298872
rect 204249 293147 204297 293175
rect 204325 293147 204359 293175
rect 204387 293147 204421 293175
rect 204449 293147 204483 293175
rect 204511 293147 204559 293175
rect 204249 293113 204559 293147
rect 204249 293085 204297 293113
rect 204325 293085 204359 293113
rect 204387 293085 204421 293113
rect 204449 293085 204483 293113
rect 204511 293085 204559 293113
rect 204249 293051 204559 293085
rect 204249 293023 204297 293051
rect 204325 293023 204359 293051
rect 204387 293023 204421 293051
rect 204449 293023 204483 293051
rect 204511 293023 204559 293051
rect 204249 292989 204559 293023
rect 204249 292961 204297 292989
rect 204325 292961 204359 292989
rect 204387 292961 204421 292989
rect 204449 292961 204483 292989
rect 204511 292961 204559 292989
rect 204249 284175 204559 292961
rect 204249 284147 204297 284175
rect 204325 284147 204359 284175
rect 204387 284147 204421 284175
rect 204449 284147 204483 284175
rect 204511 284147 204559 284175
rect 204249 284113 204559 284147
rect 204249 284085 204297 284113
rect 204325 284085 204359 284113
rect 204387 284085 204421 284113
rect 204449 284085 204483 284113
rect 204511 284085 204559 284113
rect 204249 284051 204559 284085
rect 204249 284023 204297 284051
rect 204325 284023 204359 284051
rect 204387 284023 204421 284051
rect 204449 284023 204483 284051
rect 204511 284023 204559 284051
rect 204249 283989 204559 284023
rect 204249 283961 204297 283989
rect 204325 283961 204359 283989
rect 204387 283961 204421 283989
rect 204449 283961 204483 283989
rect 204511 283961 204559 283989
rect 204249 275175 204559 283961
rect 204249 275147 204297 275175
rect 204325 275147 204359 275175
rect 204387 275147 204421 275175
rect 204449 275147 204483 275175
rect 204511 275147 204559 275175
rect 204249 275113 204559 275147
rect 204249 275085 204297 275113
rect 204325 275085 204359 275113
rect 204387 275085 204421 275113
rect 204449 275085 204483 275113
rect 204511 275085 204559 275113
rect 204249 275051 204559 275085
rect 204249 275023 204297 275051
rect 204325 275023 204359 275051
rect 204387 275023 204421 275051
rect 204449 275023 204483 275051
rect 204511 275023 204559 275051
rect 204249 274989 204559 275023
rect 204249 274961 204297 274989
rect 204325 274961 204359 274989
rect 204387 274961 204421 274989
rect 204449 274961 204483 274989
rect 204511 274961 204559 274989
rect 204249 266175 204559 274961
rect 204249 266147 204297 266175
rect 204325 266147 204359 266175
rect 204387 266147 204421 266175
rect 204449 266147 204483 266175
rect 204511 266147 204559 266175
rect 204249 266113 204559 266147
rect 204249 266085 204297 266113
rect 204325 266085 204359 266113
rect 204387 266085 204421 266113
rect 204449 266085 204483 266113
rect 204511 266085 204559 266113
rect 204249 266051 204559 266085
rect 204249 266023 204297 266051
rect 204325 266023 204359 266051
rect 204387 266023 204421 266051
rect 204449 266023 204483 266051
rect 204511 266023 204559 266051
rect 204249 265989 204559 266023
rect 204249 265961 204297 265989
rect 204325 265961 204359 265989
rect 204387 265961 204421 265989
rect 204449 265961 204483 265989
rect 204511 265961 204559 265989
rect 204249 257175 204559 265961
rect 204249 257147 204297 257175
rect 204325 257147 204359 257175
rect 204387 257147 204421 257175
rect 204449 257147 204483 257175
rect 204511 257147 204559 257175
rect 204249 257113 204559 257147
rect 204249 257085 204297 257113
rect 204325 257085 204359 257113
rect 204387 257085 204421 257113
rect 204449 257085 204483 257113
rect 204511 257085 204559 257113
rect 204249 257051 204559 257085
rect 204249 257023 204297 257051
rect 204325 257023 204359 257051
rect 204387 257023 204421 257051
rect 204449 257023 204483 257051
rect 204511 257023 204559 257051
rect 204249 256989 204559 257023
rect 204249 256961 204297 256989
rect 204325 256961 204359 256989
rect 204387 256961 204421 256989
rect 204449 256961 204483 256989
rect 204511 256961 204559 256989
rect 204249 248175 204559 256961
rect 204249 248147 204297 248175
rect 204325 248147 204359 248175
rect 204387 248147 204421 248175
rect 204449 248147 204483 248175
rect 204511 248147 204559 248175
rect 204249 248113 204559 248147
rect 204249 248085 204297 248113
rect 204325 248085 204359 248113
rect 204387 248085 204421 248113
rect 204449 248085 204483 248113
rect 204511 248085 204559 248113
rect 204249 248051 204559 248085
rect 204249 248023 204297 248051
rect 204325 248023 204359 248051
rect 204387 248023 204421 248051
rect 204449 248023 204483 248051
rect 204511 248023 204559 248051
rect 204249 247989 204559 248023
rect 204249 247961 204297 247989
rect 204325 247961 204359 247989
rect 204387 247961 204421 247989
rect 204449 247961 204483 247989
rect 204511 247961 204559 247989
rect 204249 239175 204559 247961
rect 204249 239147 204297 239175
rect 204325 239147 204359 239175
rect 204387 239147 204421 239175
rect 204449 239147 204483 239175
rect 204511 239147 204559 239175
rect 204249 239113 204559 239147
rect 204249 239085 204297 239113
rect 204325 239085 204359 239113
rect 204387 239085 204421 239113
rect 204449 239085 204483 239113
rect 204511 239085 204559 239113
rect 204249 239051 204559 239085
rect 204249 239023 204297 239051
rect 204325 239023 204359 239051
rect 204387 239023 204421 239051
rect 204449 239023 204483 239051
rect 204511 239023 204559 239051
rect 204249 238989 204559 239023
rect 204249 238961 204297 238989
rect 204325 238961 204359 238989
rect 204387 238961 204421 238989
rect 204449 238961 204483 238989
rect 204511 238961 204559 238989
rect 204249 230175 204559 238961
rect 204249 230147 204297 230175
rect 204325 230147 204359 230175
rect 204387 230147 204421 230175
rect 204449 230147 204483 230175
rect 204511 230147 204559 230175
rect 204249 230113 204559 230147
rect 204249 230085 204297 230113
rect 204325 230085 204359 230113
rect 204387 230085 204421 230113
rect 204449 230085 204483 230113
rect 204511 230085 204559 230113
rect 204249 230051 204559 230085
rect 204249 230023 204297 230051
rect 204325 230023 204359 230051
rect 204387 230023 204421 230051
rect 204449 230023 204483 230051
rect 204511 230023 204559 230051
rect 204249 229989 204559 230023
rect 204249 229961 204297 229989
rect 204325 229961 204359 229989
rect 204387 229961 204421 229989
rect 204449 229961 204483 229989
rect 204511 229961 204559 229989
rect 204249 221175 204559 229961
rect 204249 221147 204297 221175
rect 204325 221147 204359 221175
rect 204387 221147 204421 221175
rect 204449 221147 204483 221175
rect 204511 221147 204559 221175
rect 204249 221113 204559 221147
rect 204249 221085 204297 221113
rect 204325 221085 204359 221113
rect 204387 221085 204421 221113
rect 204449 221085 204483 221113
rect 204511 221085 204559 221113
rect 204249 221051 204559 221085
rect 204249 221023 204297 221051
rect 204325 221023 204359 221051
rect 204387 221023 204421 221051
rect 204449 221023 204483 221051
rect 204511 221023 204559 221051
rect 204249 220989 204559 221023
rect 204249 220961 204297 220989
rect 204325 220961 204359 220989
rect 204387 220961 204421 220989
rect 204449 220961 204483 220989
rect 204511 220961 204559 220989
rect 204249 212175 204559 220961
rect 204249 212147 204297 212175
rect 204325 212147 204359 212175
rect 204387 212147 204421 212175
rect 204449 212147 204483 212175
rect 204511 212147 204559 212175
rect 204249 212113 204559 212147
rect 204249 212085 204297 212113
rect 204325 212085 204359 212113
rect 204387 212085 204421 212113
rect 204449 212085 204483 212113
rect 204511 212085 204559 212113
rect 204249 212051 204559 212085
rect 204249 212023 204297 212051
rect 204325 212023 204359 212051
rect 204387 212023 204421 212051
rect 204449 212023 204483 212051
rect 204511 212023 204559 212051
rect 204249 211989 204559 212023
rect 204249 211961 204297 211989
rect 204325 211961 204359 211989
rect 204387 211961 204421 211989
rect 204449 211961 204483 211989
rect 204511 211961 204559 211989
rect 204249 203175 204559 211961
rect 204249 203147 204297 203175
rect 204325 203147 204359 203175
rect 204387 203147 204421 203175
rect 204449 203147 204483 203175
rect 204511 203147 204559 203175
rect 204249 203113 204559 203147
rect 204249 203085 204297 203113
rect 204325 203085 204359 203113
rect 204387 203085 204421 203113
rect 204449 203085 204483 203113
rect 204511 203085 204559 203113
rect 204249 203051 204559 203085
rect 204249 203023 204297 203051
rect 204325 203023 204359 203051
rect 204387 203023 204421 203051
rect 204449 203023 204483 203051
rect 204511 203023 204559 203051
rect 204249 202989 204559 203023
rect 204249 202961 204297 202989
rect 204325 202961 204359 202989
rect 204387 202961 204421 202989
rect 204449 202961 204483 202989
rect 204511 202961 204559 202989
rect 204249 194175 204559 202961
rect 204249 194147 204297 194175
rect 204325 194147 204359 194175
rect 204387 194147 204421 194175
rect 204449 194147 204483 194175
rect 204511 194147 204559 194175
rect 204249 194113 204559 194147
rect 204249 194085 204297 194113
rect 204325 194085 204359 194113
rect 204387 194085 204421 194113
rect 204449 194085 204483 194113
rect 204511 194085 204559 194113
rect 204249 194051 204559 194085
rect 204249 194023 204297 194051
rect 204325 194023 204359 194051
rect 204387 194023 204421 194051
rect 204449 194023 204483 194051
rect 204511 194023 204559 194051
rect 204249 193989 204559 194023
rect 204249 193961 204297 193989
rect 204325 193961 204359 193989
rect 204387 193961 204421 193989
rect 204449 193961 204483 193989
rect 204511 193961 204559 193989
rect 204249 185175 204559 193961
rect 204249 185147 204297 185175
rect 204325 185147 204359 185175
rect 204387 185147 204421 185175
rect 204449 185147 204483 185175
rect 204511 185147 204559 185175
rect 204249 185113 204559 185147
rect 204249 185085 204297 185113
rect 204325 185085 204359 185113
rect 204387 185085 204421 185113
rect 204449 185085 204483 185113
rect 204511 185085 204559 185113
rect 204249 185051 204559 185085
rect 204249 185023 204297 185051
rect 204325 185023 204359 185051
rect 204387 185023 204421 185051
rect 204449 185023 204483 185051
rect 204511 185023 204559 185051
rect 204249 184989 204559 185023
rect 204249 184961 204297 184989
rect 204325 184961 204359 184989
rect 204387 184961 204421 184989
rect 204449 184961 204483 184989
rect 204511 184961 204559 184989
rect 204249 176175 204559 184961
rect 204249 176147 204297 176175
rect 204325 176147 204359 176175
rect 204387 176147 204421 176175
rect 204449 176147 204483 176175
rect 204511 176147 204559 176175
rect 204249 176113 204559 176147
rect 204249 176085 204297 176113
rect 204325 176085 204359 176113
rect 204387 176085 204421 176113
rect 204449 176085 204483 176113
rect 204511 176085 204559 176113
rect 204249 176051 204559 176085
rect 204249 176023 204297 176051
rect 204325 176023 204359 176051
rect 204387 176023 204421 176051
rect 204449 176023 204483 176051
rect 204511 176023 204559 176051
rect 204249 175989 204559 176023
rect 204249 175961 204297 175989
rect 204325 175961 204359 175989
rect 204387 175961 204421 175989
rect 204449 175961 204483 175989
rect 204511 175961 204559 175989
rect 204249 167175 204559 175961
rect 204249 167147 204297 167175
rect 204325 167147 204359 167175
rect 204387 167147 204421 167175
rect 204449 167147 204483 167175
rect 204511 167147 204559 167175
rect 204249 167113 204559 167147
rect 204249 167085 204297 167113
rect 204325 167085 204359 167113
rect 204387 167085 204421 167113
rect 204449 167085 204483 167113
rect 204511 167085 204559 167113
rect 204249 167051 204559 167085
rect 204249 167023 204297 167051
rect 204325 167023 204359 167051
rect 204387 167023 204421 167051
rect 204449 167023 204483 167051
rect 204511 167023 204559 167051
rect 204249 166989 204559 167023
rect 204249 166961 204297 166989
rect 204325 166961 204359 166989
rect 204387 166961 204421 166989
rect 204449 166961 204483 166989
rect 204511 166961 204559 166989
rect 96729 158147 96777 158175
rect 96805 158147 96839 158175
rect 96867 158147 96901 158175
rect 96929 158147 96963 158175
rect 96991 158147 97039 158175
rect 96729 158113 97039 158147
rect 96729 158085 96777 158113
rect 96805 158085 96839 158113
rect 96867 158085 96901 158113
rect 96929 158085 96963 158113
rect 96991 158085 97039 158113
rect 96729 158051 97039 158085
rect 96729 158023 96777 158051
rect 96805 158023 96839 158051
rect 96867 158023 96901 158051
rect 96929 158023 96963 158051
rect 96991 158023 97039 158051
rect 96729 157989 97039 158023
rect 96729 157961 96777 157989
rect 96805 157961 96839 157989
rect 96867 157961 96901 157989
rect 96929 157961 96963 157989
rect 96991 157961 97039 157989
rect 96729 149175 97039 157961
rect 101344 158175 101504 158192
rect 101344 158147 101379 158175
rect 101407 158147 101441 158175
rect 101469 158147 101504 158175
rect 101344 158113 101504 158147
rect 101344 158085 101379 158113
rect 101407 158085 101441 158113
rect 101469 158085 101504 158113
rect 101344 158051 101504 158085
rect 101344 158023 101379 158051
rect 101407 158023 101441 158051
rect 101469 158023 101504 158051
rect 101344 157989 101504 158023
rect 101344 157961 101379 157989
rect 101407 157961 101441 157989
rect 101469 157961 101504 157989
rect 101344 157944 101504 157961
rect 116704 158175 116864 158192
rect 116704 158147 116739 158175
rect 116767 158147 116801 158175
rect 116829 158147 116864 158175
rect 116704 158113 116864 158147
rect 116704 158085 116739 158113
rect 116767 158085 116801 158113
rect 116829 158085 116864 158113
rect 116704 158051 116864 158085
rect 116704 158023 116739 158051
rect 116767 158023 116801 158051
rect 116829 158023 116864 158051
rect 116704 157989 116864 158023
rect 116704 157961 116739 157989
rect 116767 157961 116801 157989
rect 116829 157961 116864 157989
rect 116704 157944 116864 157961
rect 132064 158175 132224 158192
rect 132064 158147 132099 158175
rect 132127 158147 132161 158175
rect 132189 158147 132224 158175
rect 132064 158113 132224 158147
rect 132064 158085 132099 158113
rect 132127 158085 132161 158113
rect 132189 158085 132224 158113
rect 132064 158051 132224 158085
rect 132064 158023 132099 158051
rect 132127 158023 132161 158051
rect 132189 158023 132224 158051
rect 132064 157989 132224 158023
rect 132064 157961 132099 157989
rect 132127 157961 132161 157989
rect 132189 157961 132224 157989
rect 132064 157944 132224 157961
rect 147424 158175 147584 158192
rect 147424 158147 147459 158175
rect 147487 158147 147521 158175
rect 147549 158147 147584 158175
rect 147424 158113 147584 158147
rect 147424 158085 147459 158113
rect 147487 158085 147521 158113
rect 147549 158085 147584 158113
rect 147424 158051 147584 158085
rect 147424 158023 147459 158051
rect 147487 158023 147521 158051
rect 147549 158023 147584 158051
rect 147424 157989 147584 158023
rect 147424 157961 147459 157989
rect 147487 157961 147521 157989
rect 147549 157961 147584 157989
rect 147424 157944 147584 157961
rect 162784 158175 162944 158192
rect 162784 158147 162819 158175
rect 162847 158147 162881 158175
rect 162909 158147 162944 158175
rect 162784 158113 162944 158147
rect 162784 158085 162819 158113
rect 162847 158085 162881 158113
rect 162909 158085 162944 158113
rect 162784 158051 162944 158085
rect 162784 158023 162819 158051
rect 162847 158023 162881 158051
rect 162909 158023 162944 158051
rect 162784 157989 162944 158023
rect 162784 157961 162819 157989
rect 162847 157961 162881 157989
rect 162909 157961 162944 157989
rect 162784 157944 162944 157961
rect 178144 158175 178304 158192
rect 178144 158147 178179 158175
rect 178207 158147 178241 158175
rect 178269 158147 178304 158175
rect 178144 158113 178304 158147
rect 178144 158085 178179 158113
rect 178207 158085 178241 158113
rect 178269 158085 178304 158113
rect 178144 158051 178304 158085
rect 178144 158023 178179 158051
rect 178207 158023 178241 158051
rect 178269 158023 178304 158051
rect 178144 157989 178304 158023
rect 178144 157961 178179 157989
rect 178207 157961 178241 157989
rect 178269 157961 178304 157989
rect 178144 157944 178304 157961
rect 193504 158175 193664 158192
rect 193504 158147 193539 158175
rect 193567 158147 193601 158175
rect 193629 158147 193664 158175
rect 193504 158113 193664 158147
rect 193504 158085 193539 158113
rect 193567 158085 193601 158113
rect 193629 158085 193664 158113
rect 193504 158051 193664 158085
rect 193504 158023 193539 158051
rect 193567 158023 193601 158051
rect 193629 158023 193664 158051
rect 193504 157989 193664 158023
rect 193504 157961 193539 157989
rect 193567 157961 193601 157989
rect 193629 157961 193664 157989
rect 193504 157944 193664 157961
rect 204249 158175 204559 166961
rect 217749 298606 218059 299134
rect 217749 298578 217797 298606
rect 217825 298578 217859 298606
rect 217887 298578 217921 298606
rect 217949 298578 217983 298606
rect 218011 298578 218059 298606
rect 217749 298544 218059 298578
rect 217749 298516 217797 298544
rect 217825 298516 217859 298544
rect 217887 298516 217921 298544
rect 217949 298516 217983 298544
rect 218011 298516 218059 298544
rect 217749 298482 218059 298516
rect 217749 298454 217797 298482
rect 217825 298454 217859 298482
rect 217887 298454 217921 298482
rect 217949 298454 217983 298482
rect 218011 298454 218059 298482
rect 217749 298420 218059 298454
rect 217749 298392 217797 298420
rect 217825 298392 217859 298420
rect 217887 298392 217921 298420
rect 217949 298392 217983 298420
rect 218011 298392 218059 298420
rect 217749 290175 218059 298392
rect 217749 290147 217797 290175
rect 217825 290147 217859 290175
rect 217887 290147 217921 290175
rect 217949 290147 217983 290175
rect 218011 290147 218059 290175
rect 217749 290113 218059 290147
rect 217749 290085 217797 290113
rect 217825 290085 217859 290113
rect 217887 290085 217921 290113
rect 217949 290085 217983 290113
rect 218011 290085 218059 290113
rect 217749 290051 218059 290085
rect 217749 290023 217797 290051
rect 217825 290023 217859 290051
rect 217887 290023 217921 290051
rect 217949 290023 217983 290051
rect 218011 290023 218059 290051
rect 217749 289989 218059 290023
rect 217749 289961 217797 289989
rect 217825 289961 217859 289989
rect 217887 289961 217921 289989
rect 217949 289961 217983 289989
rect 218011 289961 218059 289989
rect 217749 281175 218059 289961
rect 217749 281147 217797 281175
rect 217825 281147 217859 281175
rect 217887 281147 217921 281175
rect 217949 281147 217983 281175
rect 218011 281147 218059 281175
rect 217749 281113 218059 281147
rect 217749 281085 217797 281113
rect 217825 281085 217859 281113
rect 217887 281085 217921 281113
rect 217949 281085 217983 281113
rect 218011 281085 218059 281113
rect 217749 281051 218059 281085
rect 217749 281023 217797 281051
rect 217825 281023 217859 281051
rect 217887 281023 217921 281051
rect 217949 281023 217983 281051
rect 218011 281023 218059 281051
rect 217749 280989 218059 281023
rect 217749 280961 217797 280989
rect 217825 280961 217859 280989
rect 217887 280961 217921 280989
rect 217949 280961 217983 280989
rect 218011 280961 218059 280989
rect 217749 272175 218059 280961
rect 217749 272147 217797 272175
rect 217825 272147 217859 272175
rect 217887 272147 217921 272175
rect 217949 272147 217983 272175
rect 218011 272147 218059 272175
rect 217749 272113 218059 272147
rect 217749 272085 217797 272113
rect 217825 272085 217859 272113
rect 217887 272085 217921 272113
rect 217949 272085 217983 272113
rect 218011 272085 218059 272113
rect 217749 272051 218059 272085
rect 217749 272023 217797 272051
rect 217825 272023 217859 272051
rect 217887 272023 217921 272051
rect 217949 272023 217983 272051
rect 218011 272023 218059 272051
rect 217749 271989 218059 272023
rect 217749 271961 217797 271989
rect 217825 271961 217859 271989
rect 217887 271961 217921 271989
rect 217949 271961 217983 271989
rect 218011 271961 218059 271989
rect 217749 263175 218059 271961
rect 217749 263147 217797 263175
rect 217825 263147 217859 263175
rect 217887 263147 217921 263175
rect 217949 263147 217983 263175
rect 218011 263147 218059 263175
rect 217749 263113 218059 263147
rect 217749 263085 217797 263113
rect 217825 263085 217859 263113
rect 217887 263085 217921 263113
rect 217949 263085 217983 263113
rect 218011 263085 218059 263113
rect 217749 263051 218059 263085
rect 217749 263023 217797 263051
rect 217825 263023 217859 263051
rect 217887 263023 217921 263051
rect 217949 263023 217983 263051
rect 218011 263023 218059 263051
rect 217749 262989 218059 263023
rect 217749 262961 217797 262989
rect 217825 262961 217859 262989
rect 217887 262961 217921 262989
rect 217949 262961 217983 262989
rect 218011 262961 218059 262989
rect 217749 254175 218059 262961
rect 217749 254147 217797 254175
rect 217825 254147 217859 254175
rect 217887 254147 217921 254175
rect 217949 254147 217983 254175
rect 218011 254147 218059 254175
rect 217749 254113 218059 254147
rect 217749 254085 217797 254113
rect 217825 254085 217859 254113
rect 217887 254085 217921 254113
rect 217949 254085 217983 254113
rect 218011 254085 218059 254113
rect 217749 254051 218059 254085
rect 217749 254023 217797 254051
rect 217825 254023 217859 254051
rect 217887 254023 217921 254051
rect 217949 254023 217983 254051
rect 218011 254023 218059 254051
rect 217749 253989 218059 254023
rect 217749 253961 217797 253989
rect 217825 253961 217859 253989
rect 217887 253961 217921 253989
rect 217949 253961 217983 253989
rect 218011 253961 218059 253989
rect 217749 245175 218059 253961
rect 217749 245147 217797 245175
rect 217825 245147 217859 245175
rect 217887 245147 217921 245175
rect 217949 245147 217983 245175
rect 218011 245147 218059 245175
rect 217749 245113 218059 245147
rect 217749 245085 217797 245113
rect 217825 245085 217859 245113
rect 217887 245085 217921 245113
rect 217949 245085 217983 245113
rect 218011 245085 218059 245113
rect 217749 245051 218059 245085
rect 217749 245023 217797 245051
rect 217825 245023 217859 245051
rect 217887 245023 217921 245051
rect 217949 245023 217983 245051
rect 218011 245023 218059 245051
rect 217749 244989 218059 245023
rect 217749 244961 217797 244989
rect 217825 244961 217859 244989
rect 217887 244961 217921 244989
rect 217949 244961 217983 244989
rect 218011 244961 218059 244989
rect 217749 236175 218059 244961
rect 217749 236147 217797 236175
rect 217825 236147 217859 236175
rect 217887 236147 217921 236175
rect 217949 236147 217983 236175
rect 218011 236147 218059 236175
rect 217749 236113 218059 236147
rect 217749 236085 217797 236113
rect 217825 236085 217859 236113
rect 217887 236085 217921 236113
rect 217949 236085 217983 236113
rect 218011 236085 218059 236113
rect 217749 236051 218059 236085
rect 217749 236023 217797 236051
rect 217825 236023 217859 236051
rect 217887 236023 217921 236051
rect 217949 236023 217983 236051
rect 218011 236023 218059 236051
rect 217749 235989 218059 236023
rect 217749 235961 217797 235989
rect 217825 235961 217859 235989
rect 217887 235961 217921 235989
rect 217949 235961 217983 235989
rect 218011 235961 218059 235989
rect 217749 227175 218059 235961
rect 217749 227147 217797 227175
rect 217825 227147 217859 227175
rect 217887 227147 217921 227175
rect 217949 227147 217983 227175
rect 218011 227147 218059 227175
rect 217749 227113 218059 227147
rect 217749 227085 217797 227113
rect 217825 227085 217859 227113
rect 217887 227085 217921 227113
rect 217949 227085 217983 227113
rect 218011 227085 218059 227113
rect 217749 227051 218059 227085
rect 217749 227023 217797 227051
rect 217825 227023 217859 227051
rect 217887 227023 217921 227051
rect 217949 227023 217983 227051
rect 218011 227023 218059 227051
rect 217749 226989 218059 227023
rect 217749 226961 217797 226989
rect 217825 226961 217859 226989
rect 217887 226961 217921 226989
rect 217949 226961 217983 226989
rect 218011 226961 218059 226989
rect 217749 218175 218059 226961
rect 217749 218147 217797 218175
rect 217825 218147 217859 218175
rect 217887 218147 217921 218175
rect 217949 218147 217983 218175
rect 218011 218147 218059 218175
rect 217749 218113 218059 218147
rect 217749 218085 217797 218113
rect 217825 218085 217859 218113
rect 217887 218085 217921 218113
rect 217949 218085 217983 218113
rect 218011 218085 218059 218113
rect 217749 218051 218059 218085
rect 217749 218023 217797 218051
rect 217825 218023 217859 218051
rect 217887 218023 217921 218051
rect 217949 218023 217983 218051
rect 218011 218023 218059 218051
rect 217749 217989 218059 218023
rect 217749 217961 217797 217989
rect 217825 217961 217859 217989
rect 217887 217961 217921 217989
rect 217949 217961 217983 217989
rect 218011 217961 218059 217989
rect 217749 209175 218059 217961
rect 217749 209147 217797 209175
rect 217825 209147 217859 209175
rect 217887 209147 217921 209175
rect 217949 209147 217983 209175
rect 218011 209147 218059 209175
rect 217749 209113 218059 209147
rect 217749 209085 217797 209113
rect 217825 209085 217859 209113
rect 217887 209085 217921 209113
rect 217949 209085 217983 209113
rect 218011 209085 218059 209113
rect 217749 209051 218059 209085
rect 217749 209023 217797 209051
rect 217825 209023 217859 209051
rect 217887 209023 217921 209051
rect 217949 209023 217983 209051
rect 218011 209023 218059 209051
rect 217749 208989 218059 209023
rect 217749 208961 217797 208989
rect 217825 208961 217859 208989
rect 217887 208961 217921 208989
rect 217949 208961 217983 208989
rect 218011 208961 218059 208989
rect 217749 200175 218059 208961
rect 217749 200147 217797 200175
rect 217825 200147 217859 200175
rect 217887 200147 217921 200175
rect 217949 200147 217983 200175
rect 218011 200147 218059 200175
rect 217749 200113 218059 200147
rect 217749 200085 217797 200113
rect 217825 200085 217859 200113
rect 217887 200085 217921 200113
rect 217949 200085 217983 200113
rect 218011 200085 218059 200113
rect 217749 200051 218059 200085
rect 217749 200023 217797 200051
rect 217825 200023 217859 200051
rect 217887 200023 217921 200051
rect 217949 200023 217983 200051
rect 218011 200023 218059 200051
rect 217749 199989 218059 200023
rect 217749 199961 217797 199989
rect 217825 199961 217859 199989
rect 217887 199961 217921 199989
rect 217949 199961 217983 199989
rect 218011 199961 218059 199989
rect 217749 191175 218059 199961
rect 217749 191147 217797 191175
rect 217825 191147 217859 191175
rect 217887 191147 217921 191175
rect 217949 191147 217983 191175
rect 218011 191147 218059 191175
rect 217749 191113 218059 191147
rect 217749 191085 217797 191113
rect 217825 191085 217859 191113
rect 217887 191085 217921 191113
rect 217949 191085 217983 191113
rect 218011 191085 218059 191113
rect 217749 191051 218059 191085
rect 217749 191023 217797 191051
rect 217825 191023 217859 191051
rect 217887 191023 217921 191051
rect 217949 191023 217983 191051
rect 218011 191023 218059 191051
rect 217749 190989 218059 191023
rect 217749 190961 217797 190989
rect 217825 190961 217859 190989
rect 217887 190961 217921 190989
rect 217949 190961 217983 190989
rect 218011 190961 218059 190989
rect 217749 182175 218059 190961
rect 217749 182147 217797 182175
rect 217825 182147 217859 182175
rect 217887 182147 217921 182175
rect 217949 182147 217983 182175
rect 218011 182147 218059 182175
rect 217749 182113 218059 182147
rect 217749 182085 217797 182113
rect 217825 182085 217859 182113
rect 217887 182085 217921 182113
rect 217949 182085 217983 182113
rect 218011 182085 218059 182113
rect 217749 182051 218059 182085
rect 217749 182023 217797 182051
rect 217825 182023 217859 182051
rect 217887 182023 217921 182051
rect 217949 182023 217983 182051
rect 218011 182023 218059 182051
rect 217749 181989 218059 182023
rect 217749 181961 217797 181989
rect 217825 181961 217859 181989
rect 217887 181961 217921 181989
rect 217949 181961 217983 181989
rect 218011 181961 218059 181989
rect 217749 173175 218059 181961
rect 217749 173147 217797 173175
rect 217825 173147 217859 173175
rect 217887 173147 217921 173175
rect 217949 173147 217983 173175
rect 218011 173147 218059 173175
rect 217749 173113 218059 173147
rect 217749 173085 217797 173113
rect 217825 173085 217859 173113
rect 217887 173085 217921 173113
rect 217949 173085 217983 173113
rect 218011 173085 218059 173113
rect 217749 173051 218059 173085
rect 217749 173023 217797 173051
rect 217825 173023 217859 173051
rect 217887 173023 217921 173051
rect 217949 173023 217983 173051
rect 218011 173023 218059 173051
rect 217749 172989 218059 173023
rect 217749 172961 217797 172989
rect 217825 172961 217859 172989
rect 217887 172961 217921 172989
rect 217949 172961 217983 172989
rect 218011 172961 218059 172989
rect 217749 164175 218059 172961
rect 217749 164147 217797 164175
rect 217825 164147 217859 164175
rect 217887 164147 217921 164175
rect 217949 164147 217983 164175
rect 218011 164147 218059 164175
rect 217749 164113 218059 164147
rect 217749 164085 217797 164113
rect 217825 164085 217859 164113
rect 217887 164085 217921 164113
rect 217949 164085 217983 164113
rect 218011 164085 218059 164113
rect 217749 164051 218059 164085
rect 217749 164023 217797 164051
rect 217825 164023 217859 164051
rect 217887 164023 217921 164051
rect 217949 164023 217983 164051
rect 218011 164023 218059 164051
rect 217749 163989 218059 164023
rect 217749 163961 217797 163989
rect 217825 163961 217859 163989
rect 217887 163961 217921 163989
rect 217949 163961 217983 163989
rect 218011 163961 218059 163989
rect 207046 162050 207074 162055
rect 207046 161770 207074 162022
rect 207046 161737 207074 161742
rect 204249 158147 204297 158175
rect 204325 158147 204359 158175
rect 204387 158147 204421 158175
rect 204449 158147 204483 158175
rect 204511 158147 204559 158175
rect 204249 158113 204559 158147
rect 204249 158085 204297 158113
rect 204325 158085 204359 158113
rect 204387 158085 204421 158113
rect 204449 158085 204483 158113
rect 204511 158085 204559 158113
rect 204249 158051 204559 158085
rect 204249 158023 204297 158051
rect 204325 158023 204359 158051
rect 204387 158023 204421 158051
rect 204449 158023 204483 158051
rect 204511 158023 204559 158051
rect 204249 157989 204559 158023
rect 204249 157961 204297 157989
rect 204325 157961 204359 157989
rect 204387 157961 204421 157989
rect 204449 157961 204483 157989
rect 204511 157961 204559 157989
rect 109024 155175 109184 155192
rect 109024 155147 109059 155175
rect 109087 155147 109121 155175
rect 109149 155147 109184 155175
rect 109024 155113 109184 155147
rect 109024 155085 109059 155113
rect 109087 155085 109121 155113
rect 109149 155085 109184 155113
rect 109024 155051 109184 155085
rect 109024 155023 109059 155051
rect 109087 155023 109121 155051
rect 109149 155023 109184 155051
rect 109024 154989 109184 155023
rect 109024 154961 109059 154989
rect 109087 154961 109121 154989
rect 109149 154961 109184 154989
rect 109024 154944 109184 154961
rect 124384 155175 124544 155192
rect 124384 155147 124419 155175
rect 124447 155147 124481 155175
rect 124509 155147 124544 155175
rect 124384 155113 124544 155147
rect 124384 155085 124419 155113
rect 124447 155085 124481 155113
rect 124509 155085 124544 155113
rect 124384 155051 124544 155085
rect 124384 155023 124419 155051
rect 124447 155023 124481 155051
rect 124509 155023 124544 155051
rect 124384 154989 124544 155023
rect 124384 154961 124419 154989
rect 124447 154961 124481 154989
rect 124509 154961 124544 154989
rect 124384 154944 124544 154961
rect 139744 155175 139904 155192
rect 139744 155147 139779 155175
rect 139807 155147 139841 155175
rect 139869 155147 139904 155175
rect 139744 155113 139904 155147
rect 139744 155085 139779 155113
rect 139807 155085 139841 155113
rect 139869 155085 139904 155113
rect 139744 155051 139904 155085
rect 139744 155023 139779 155051
rect 139807 155023 139841 155051
rect 139869 155023 139904 155051
rect 139744 154989 139904 155023
rect 139744 154961 139779 154989
rect 139807 154961 139841 154989
rect 139869 154961 139904 154989
rect 139744 154944 139904 154961
rect 155104 155175 155264 155192
rect 155104 155147 155139 155175
rect 155167 155147 155201 155175
rect 155229 155147 155264 155175
rect 155104 155113 155264 155147
rect 155104 155085 155139 155113
rect 155167 155085 155201 155113
rect 155229 155085 155264 155113
rect 155104 155051 155264 155085
rect 155104 155023 155139 155051
rect 155167 155023 155201 155051
rect 155229 155023 155264 155051
rect 155104 154989 155264 155023
rect 155104 154961 155139 154989
rect 155167 154961 155201 154989
rect 155229 154961 155264 154989
rect 155104 154944 155264 154961
rect 170464 155175 170624 155192
rect 170464 155147 170499 155175
rect 170527 155147 170561 155175
rect 170589 155147 170624 155175
rect 170464 155113 170624 155147
rect 170464 155085 170499 155113
rect 170527 155085 170561 155113
rect 170589 155085 170624 155113
rect 170464 155051 170624 155085
rect 170464 155023 170499 155051
rect 170527 155023 170561 155051
rect 170589 155023 170624 155051
rect 170464 154989 170624 155023
rect 170464 154961 170499 154989
rect 170527 154961 170561 154989
rect 170589 154961 170624 154989
rect 170464 154944 170624 154961
rect 185824 155175 185984 155192
rect 185824 155147 185859 155175
rect 185887 155147 185921 155175
rect 185949 155147 185984 155175
rect 185824 155113 185984 155147
rect 185824 155085 185859 155113
rect 185887 155085 185921 155113
rect 185949 155085 185984 155113
rect 185824 155051 185984 155085
rect 185824 155023 185859 155051
rect 185887 155023 185921 155051
rect 185949 155023 185984 155051
rect 185824 154989 185984 155023
rect 185824 154961 185859 154989
rect 185887 154961 185921 154989
rect 185949 154961 185984 154989
rect 185824 154944 185984 154961
rect 201184 155175 201344 155192
rect 201184 155147 201219 155175
rect 201247 155147 201281 155175
rect 201309 155147 201344 155175
rect 201184 155113 201344 155147
rect 201184 155085 201219 155113
rect 201247 155085 201281 155113
rect 201309 155085 201344 155113
rect 201184 155051 201344 155085
rect 201184 155023 201219 155051
rect 201247 155023 201281 155051
rect 201309 155023 201344 155051
rect 201184 154989 201344 155023
rect 201184 154961 201219 154989
rect 201247 154961 201281 154989
rect 201309 154961 201344 154989
rect 201184 154944 201344 154961
rect 96729 149147 96777 149175
rect 96805 149147 96839 149175
rect 96867 149147 96901 149175
rect 96929 149147 96963 149175
rect 96991 149147 97039 149175
rect 96729 149113 97039 149147
rect 96729 149085 96777 149113
rect 96805 149085 96839 149113
rect 96867 149085 96901 149113
rect 96929 149085 96963 149113
rect 96991 149085 97039 149113
rect 96729 149051 97039 149085
rect 96729 149023 96777 149051
rect 96805 149023 96839 149051
rect 96867 149023 96901 149051
rect 96929 149023 96963 149051
rect 96991 149023 97039 149051
rect 96729 148989 97039 149023
rect 96729 148961 96777 148989
rect 96805 148961 96839 148989
rect 96867 148961 96901 148989
rect 96929 148961 96963 148989
rect 96991 148961 97039 148989
rect 96729 140175 97039 148961
rect 101344 149175 101504 149192
rect 101344 149147 101379 149175
rect 101407 149147 101441 149175
rect 101469 149147 101504 149175
rect 101344 149113 101504 149147
rect 101344 149085 101379 149113
rect 101407 149085 101441 149113
rect 101469 149085 101504 149113
rect 101344 149051 101504 149085
rect 101344 149023 101379 149051
rect 101407 149023 101441 149051
rect 101469 149023 101504 149051
rect 101344 148989 101504 149023
rect 101344 148961 101379 148989
rect 101407 148961 101441 148989
rect 101469 148961 101504 148989
rect 101344 148944 101504 148961
rect 116704 149175 116864 149192
rect 116704 149147 116739 149175
rect 116767 149147 116801 149175
rect 116829 149147 116864 149175
rect 116704 149113 116864 149147
rect 116704 149085 116739 149113
rect 116767 149085 116801 149113
rect 116829 149085 116864 149113
rect 116704 149051 116864 149085
rect 116704 149023 116739 149051
rect 116767 149023 116801 149051
rect 116829 149023 116864 149051
rect 116704 148989 116864 149023
rect 116704 148961 116739 148989
rect 116767 148961 116801 148989
rect 116829 148961 116864 148989
rect 116704 148944 116864 148961
rect 132064 149175 132224 149192
rect 132064 149147 132099 149175
rect 132127 149147 132161 149175
rect 132189 149147 132224 149175
rect 132064 149113 132224 149147
rect 132064 149085 132099 149113
rect 132127 149085 132161 149113
rect 132189 149085 132224 149113
rect 132064 149051 132224 149085
rect 132064 149023 132099 149051
rect 132127 149023 132161 149051
rect 132189 149023 132224 149051
rect 132064 148989 132224 149023
rect 132064 148961 132099 148989
rect 132127 148961 132161 148989
rect 132189 148961 132224 148989
rect 132064 148944 132224 148961
rect 147424 149175 147584 149192
rect 147424 149147 147459 149175
rect 147487 149147 147521 149175
rect 147549 149147 147584 149175
rect 147424 149113 147584 149147
rect 147424 149085 147459 149113
rect 147487 149085 147521 149113
rect 147549 149085 147584 149113
rect 147424 149051 147584 149085
rect 147424 149023 147459 149051
rect 147487 149023 147521 149051
rect 147549 149023 147584 149051
rect 147424 148989 147584 149023
rect 147424 148961 147459 148989
rect 147487 148961 147521 148989
rect 147549 148961 147584 148989
rect 147424 148944 147584 148961
rect 162784 149175 162944 149192
rect 162784 149147 162819 149175
rect 162847 149147 162881 149175
rect 162909 149147 162944 149175
rect 162784 149113 162944 149147
rect 162784 149085 162819 149113
rect 162847 149085 162881 149113
rect 162909 149085 162944 149113
rect 162784 149051 162944 149085
rect 162784 149023 162819 149051
rect 162847 149023 162881 149051
rect 162909 149023 162944 149051
rect 162784 148989 162944 149023
rect 162784 148961 162819 148989
rect 162847 148961 162881 148989
rect 162909 148961 162944 148989
rect 162784 148944 162944 148961
rect 178144 149175 178304 149192
rect 178144 149147 178179 149175
rect 178207 149147 178241 149175
rect 178269 149147 178304 149175
rect 178144 149113 178304 149147
rect 178144 149085 178179 149113
rect 178207 149085 178241 149113
rect 178269 149085 178304 149113
rect 178144 149051 178304 149085
rect 178144 149023 178179 149051
rect 178207 149023 178241 149051
rect 178269 149023 178304 149051
rect 178144 148989 178304 149023
rect 178144 148961 178179 148989
rect 178207 148961 178241 148989
rect 178269 148961 178304 148989
rect 178144 148944 178304 148961
rect 193504 149175 193664 149192
rect 193504 149147 193539 149175
rect 193567 149147 193601 149175
rect 193629 149147 193664 149175
rect 193504 149113 193664 149147
rect 193504 149085 193539 149113
rect 193567 149085 193601 149113
rect 193629 149085 193664 149113
rect 193504 149051 193664 149085
rect 193504 149023 193539 149051
rect 193567 149023 193601 149051
rect 193629 149023 193664 149051
rect 193504 148989 193664 149023
rect 193504 148961 193539 148989
rect 193567 148961 193601 148989
rect 193629 148961 193664 148989
rect 193504 148944 193664 148961
rect 204249 149175 204559 157961
rect 208864 158175 209024 158192
rect 208864 158147 208899 158175
rect 208927 158147 208961 158175
rect 208989 158147 209024 158175
rect 208864 158113 209024 158147
rect 208864 158085 208899 158113
rect 208927 158085 208961 158113
rect 208989 158085 209024 158113
rect 208864 158051 209024 158085
rect 208864 158023 208899 158051
rect 208927 158023 208961 158051
rect 208989 158023 209024 158051
rect 208864 157989 209024 158023
rect 208864 157961 208899 157989
rect 208927 157961 208961 157989
rect 208989 157961 209024 157989
rect 208864 157944 209024 157961
rect 216544 155175 216704 155192
rect 216544 155147 216579 155175
rect 216607 155147 216641 155175
rect 216669 155147 216704 155175
rect 216544 155113 216704 155147
rect 216544 155085 216579 155113
rect 216607 155085 216641 155113
rect 216669 155085 216704 155113
rect 216544 155051 216704 155085
rect 216544 155023 216579 155051
rect 216607 155023 216641 155051
rect 216669 155023 216704 155051
rect 216544 154989 216704 155023
rect 216544 154961 216579 154989
rect 216607 154961 216641 154989
rect 216669 154961 216704 154989
rect 216544 154944 216704 154961
rect 217749 155175 218059 163961
rect 217749 155147 217797 155175
rect 217825 155147 217859 155175
rect 217887 155147 217921 155175
rect 217949 155147 217983 155175
rect 218011 155147 218059 155175
rect 217749 155113 218059 155147
rect 217749 155085 217797 155113
rect 217825 155085 217859 155113
rect 217887 155085 217921 155113
rect 217949 155085 217983 155113
rect 218011 155085 218059 155113
rect 217749 155051 218059 155085
rect 217749 155023 217797 155051
rect 217825 155023 217859 155051
rect 217887 155023 217921 155051
rect 217949 155023 217983 155051
rect 218011 155023 218059 155051
rect 217749 154989 218059 155023
rect 217749 154961 217797 154989
rect 217825 154961 217859 154989
rect 217887 154961 217921 154989
rect 217949 154961 217983 154989
rect 218011 154961 218059 154989
rect 204249 149147 204297 149175
rect 204325 149147 204359 149175
rect 204387 149147 204421 149175
rect 204449 149147 204483 149175
rect 204511 149147 204559 149175
rect 204249 149113 204559 149147
rect 204249 149085 204297 149113
rect 204325 149085 204359 149113
rect 204387 149085 204421 149113
rect 204449 149085 204483 149113
rect 204511 149085 204559 149113
rect 204249 149051 204559 149085
rect 204249 149023 204297 149051
rect 204325 149023 204359 149051
rect 204387 149023 204421 149051
rect 204449 149023 204483 149051
rect 204511 149023 204559 149051
rect 204249 148989 204559 149023
rect 204249 148961 204297 148989
rect 204325 148961 204359 148989
rect 204387 148961 204421 148989
rect 204449 148961 204483 148989
rect 204511 148961 204559 148989
rect 109024 146175 109184 146192
rect 109024 146147 109059 146175
rect 109087 146147 109121 146175
rect 109149 146147 109184 146175
rect 109024 146113 109184 146147
rect 109024 146085 109059 146113
rect 109087 146085 109121 146113
rect 109149 146085 109184 146113
rect 109024 146051 109184 146085
rect 109024 146023 109059 146051
rect 109087 146023 109121 146051
rect 109149 146023 109184 146051
rect 109024 145989 109184 146023
rect 109024 145961 109059 145989
rect 109087 145961 109121 145989
rect 109149 145961 109184 145989
rect 109024 145944 109184 145961
rect 124384 146175 124544 146192
rect 124384 146147 124419 146175
rect 124447 146147 124481 146175
rect 124509 146147 124544 146175
rect 124384 146113 124544 146147
rect 124384 146085 124419 146113
rect 124447 146085 124481 146113
rect 124509 146085 124544 146113
rect 124384 146051 124544 146085
rect 124384 146023 124419 146051
rect 124447 146023 124481 146051
rect 124509 146023 124544 146051
rect 124384 145989 124544 146023
rect 124384 145961 124419 145989
rect 124447 145961 124481 145989
rect 124509 145961 124544 145989
rect 124384 145944 124544 145961
rect 139744 146175 139904 146192
rect 139744 146147 139779 146175
rect 139807 146147 139841 146175
rect 139869 146147 139904 146175
rect 139744 146113 139904 146147
rect 139744 146085 139779 146113
rect 139807 146085 139841 146113
rect 139869 146085 139904 146113
rect 139744 146051 139904 146085
rect 139744 146023 139779 146051
rect 139807 146023 139841 146051
rect 139869 146023 139904 146051
rect 139744 145989 139904 146023
rect 139744 145961 139779 145989
rect 139807 145961 139841 145989
rect 139869 145961 139904 145989
rect 139744 145944 139904 145961
rect 155104 146175 155264 146192
rect 155104 146147 155139 146175
rect 155167 146147 155201 146175
rect 155229 146147 155264 146175
rect 155104 146113 155264 146147
rect 155104 146085 155139 146113
rect 155167 146085 155201 146113
rect 155229 146085 155264 146113
rect 155104 146051 155264 146085
rect 155104 146023 155139 146051
rect 155167 146023 155201 146051
rect 155229 146023 155264 146051
rect 155104 145989 155264 146023
rect 155104 145961 155139 145989
rect 155167 145961 155201 145989
rect 155229 145961 155264 145989
rect 155104 145944 155264 145961
rect 170464 146175 170624 146192
rect 170464 146147 170499 146175
rect 170527 146147 170561 146175
rect 170589 146147 170624 146175
rect 170464 146113 170624 146147
rect 170464 146085 170499 146113
rect 170527 146085 170561 146113
rect 170589 146085 170624 146113
rect 170464 146051 170624 146085
rect 170464 146023 170499 146051
rect 170527 146023 170561 146051
rect 170589 146023 170624 146051
rect 170464 145989 170624 146023
rect 170464 145961 170499 145989
rect 170527 145961 170561 145989
rect 170589 145961 170624 145989
rect 170464 145944 170624 145961
rect 185824 146175 185984 146192
rect 185824 146147 185859 146175
rect 185887 146147 185921 146175
rect 185949 146147 185984 146175
rect 185824 146113 185984 146147
rect 185824 146085 185859 146113
rect 185887 146085 185921 146113
rect 185949 146085 185984 146113
rect 185824 146051 185984 146085
rect 185824 146023 185859 146051
rect 185887 146023 185921 146051
rect 185949 146023 185984 146051
rect 185824 145989 185984 146023
rect 185824 145961 185859 145989
rect 185887 145961 185921 145989
rect 185949 145961 185984 145989
rect 185824 145944 185984 145961
rect 201184 146175 201344 146192
rect 201184 146147 201219 146175
rect 201247 146147 201281 146175
rect 201309 146147 201344 146175
rect 201184 146113 201344 146147
rect 201184 146085 201219 146113
rect 201247 146085 201281 146113
rect 201309 146085 201344 146113
rect 201184 146051 201344 146085
rect 201184 146023 201219 146051
rect 201247 146023 201281 146051
rect 201309 146023 201344 146051
rect 201184 145989 201344 146023
rect 201184 145961 201219 145989
rect 201247 145961 201281 145989
rect 201309 145961 201344 145989
rect 201184 145944 201344 145961
rect 96729 140147 96777 140175
rect 96805 140147 96839 140175
rect 96867 140147 96901 140175
rect 96929 140147 96963 140175
rect 96991 140147 97039 140175
rect 96729 140113 97039 140147
rect 96729 140085 96777 140113
rect 96805 140085 96839 140113
rect 96867 140085 96901 140113
rect 96929 140085 96963 140113
rect 96991 140085 97039 140113
rect 96729 140051 97039 140085
rect 96729 140023 96777 140051
rect 96805 140023 96839 140051
rect 96867 140023 96901 140051
rect 96929 140023 96963 140051
rect 96991 140023 97039 140051
rect 96729 139989 97039 140023
rect 96729 139961 96777 139989
rect 96805 139961 96839 139989
rect 96867 139961 96901 139989
rect 96929 139961 96963 139989
rect 96991 139961 97039 139989
rect 96729 131175 97039 139961
rect 101344 140175 101504 140192
rect 101344 140147 101379 140175
rect 101407 140147 101441 140175
rect 101469 140147 101504 140175
rect 101344 140113 101504 140147
rect 101344 140085 101379 140113
rect 101407 140085 101441 140113
rect 101469 140085 101504 140113
rect 101344 140051 101504 140085
rect 101344 140023 101379 140051
rect 101407 140023 101441 140051
rect 101469 140023 101504 140051
rect 101344 139989 101504 140023
rect 101344 139961 101379 139989
rect 101407 139961 101441 139989
rect 101469 139961 101504 139989
rect 101344 139944 101504 139961
rect 116704 140175 116864 140192
rect 116704 140147 116739 140175
rect 116767 140147 116801 140175
rect 116829 140147 116864 140175
rect 116704 140113 116864 140147
rect 116704 140085 116739 140113
rect 116767 140085 116801 140113
rect 116829 140085 116864 140113
rect 116704 140051 116864 140085
rect 116704 140023 116739 140051
rect 116767 140023 116801 140051
rect 116829 140023 116864 140051
rect 116704 139989 116864 140023
rect 116704 139961 116739 139989
rect 116767 139961 116801 139989
rect 116829 139961 116864 139989
rect 116704 139944 116864 139961
rect 132064 140175 132224 140192
rect 132064 140147 132099 140175
rect 132127 140147 132161 140175
rect 132189 140147 132224 140175
rect 132064 140113 132224 140147
rect 132064 140085 132099 140113
rect 132127 140085 132161 140113
rect 132189 140085 132224 140113
rect 132064 140051 132224 140085
rect 132064 140023 132099 140051
rect 132127 140023 132161 140051
rect 132189 140023 132224 140051
rect 132064 139989 132224 140023
rect 132064 139961 132099 139989
rect 132127 139961 132161 139989
rect 132189 139961 132224 139989
rect 132064 139944 132224 139961
rect 147424 140175 147584 140192
rect 147424 140147 147459 140175
rect 147487 140147 147521 140175
rect 147549 140147 147584 140175
rect 147424 140113 147584 140147
rect 147424 140085 147459 140113
rect 147487 140085 147521 140113
rect 147549 140085 147584 140113
rect 147424 140051 147584 140085
rect 147424 140023 147459 140051
rect 147487 140023 147521 140051
rect 147549 140023 147584 140051
rect 147424 139989 147584 140023
rect 147424 139961 147459 139989
rect 147487 139961 147521 139989
rect 147549 139961 147584 139989
rect 147424 139944 147584 139961
rect 162784 140175 162944 140192
rect 162784 140147 162819 140175
rect 162847 140147 162881 140175
rect 162909 140147 162944 140175
rect 162784 140113 162944 140147
rect 162784 140085 162819 140113
rect 162847 140085 162881 140113
rect 162909 140085 162944 140113
rect 162784 140051 162944 140085
rect 162784 140023 162819 140051
rect 162847 140023 162881 140051
rect 162909 140023 162944 140051
rect 162784 139989 162944 140023
rect 162784 139961 162819 139989
rect 162847 139961 162881 139989
rect 162909 139961 162944 139989
rect 162784 139944 162944 139961
rect 178144 140175 178304 140192
rect 178144 140147 178179 140175
rect 178207 140147 178241 140175
rect 178269 140147 178304 140175
rect 178144 140113 178304 140147
rect 178144 140085 178179 140113
rect 178207 140085 178241 140113
rect 178269 140085 178304 140113
rect 178144 140051 178304 140085
rect 178144 140023 178179 140051
rect 178207 140023 178241 140051
rect 178269 140023 178304 140051
rect 178144 139989 178304 140023
rect 178144 139961 178179 139989
rect 178207 139961 178241 139989
rect 178269 139961 178304 139989
rect 178144 139944 178304 139961
rect 193504 140175 193664 140192
rect 193504 140147 193539 140175
rect 193567 140147 193601 140175
rect 193629 140147 193664 140175
rect 193504 140113 193664 140147
rect 193504 140085 193539 140113
rect 193567 140085 193601 140113
rect 193629 140085 193664 140113
rect 193504 140051 193664 140085
rect 193504 140023 193539 140051
rect 193567 140023 193601 140051
rect 193629 140023 193664 140051
rect 193504 139989 193664 140023
rect 193504 139961 193539 139989
rect 193567 139961 193601 139989
rect 193629 139961 193664 139989
rect 193504 139944 193664 139961
rect 204249 140175 204559 148961
rect 208864 149175 209024 149192
rect 208864 149147 208899 149175
rect 208927 149147 208961 149175
rect 208989 149147 209024 149175
rect 208864 149113 209024 149147
rect 208864 149085 208899 149113
rect 208927 149085 208961 149113
rect 208989 149085 209024 149113
rect 208864 149051 209024 149085
rect 208864 149023 208899 149051
rect 208927 149023 208961 149051
rect 208989 149023 209024 149051
rect 208864 148989 209024 149023
rect 208864 148961 208899 148989
rect 208927 148961 208961 148989
rect 208989 148961 209024 148989
rect 208864 148944 209024 148961
rect 216544 146175 216704 146192
rect 216544 146147 216579 146175
rect 216607 146147 216641 146175
rect 216669 146147 216704 146175
rect 216544 146113 216704 146147
rect 216544 146085 216579 146113
rect 216607 146085 216641 146113
rect 216669 146085 216704 146113
rect 216544 146051 216704 146085
rect 216544 146023 216579 146051
rect 216607 146023 216641 146051
rect 216669 146023 216704 146051
rect 216544 145989 216704 146023
rect 216544 145961 216579 145989
rect 216607 145961 216641 145989
rect 216669 145961 216704 145989
rect 216544 145944 216704 145961
rect 217749 146175 218059 154961
rect 217749 146147 217797 146175
rect 217825 146147 217859 146175
rect 217887 146147 217921 146175
rect 217949 146147 217983 146175
rect 218011 146147 218059 146175
rect 217749 146113 218059 146147
rect 217749 146085 217797 146113
rect 217825 146085 217859 146113
rect 217887 146085 217921 146113
rect 217949 146085 217983 146113
rect 218011 146085 218059 146113
rect 217749 146051 218059 146085
rect 217749 146023 217797 146051
rect 217825 146023 217859 146051
rect 217887 146023 217921 146051
rect 217949 146023 217983 146051
rect 218011 146023 218059 146051
rect 217749 145989 218059 146023
rect 217749 145961 217797 145989
rect 217825 145961 217859 145989
rect 217887 145961 217921 145989
rect 217949 145961 217983 145989
rect 218011 145961 218059 145989
rect 204249 140147 204297 140175
rect 204325 140147 204359 140175
rect 204387 140147 204421 140175
rect 204449 140147 204483 140175
rect 204511 140147 204559 140175
rect 204249 140113 204559 140147
rect 204249 140085 204297 140113
rect 204325 140085 204359 140113
rect 204387 140085 204421 140113
rect 204449 140085 204483 140113
rect 204511 140085 204559 140113
rect 204249 140051 204559 140085
rect 204249 140023 204297 140051
rect 204325 140023 204359 140051
rect 204387 140023 204421 140051
rect 204449 140023 204483 140051
rect 204511 140023 204559 140051
rect 204249 139989 204559 140023
rect 204249 139961 204297 139989
rect 204325 139961 204359 139989
rect 204387 139961 204421 139989
rect 204449 139961 204483 139989
rect 204511 139961 204559 139989
rect 109024 137175 109184 137192
rect 109024 137147 109059 137175
rect 109087 137147 109121 137175
rect 109149 137147 109184 137175
rect 109024 137113 109184 137147
rect 109024 137085 109059 137113
rect 109087 137085 109121 137113
rect 109149 137085 109184 137113
rect 109024 137051 109184 137085
rect 109024 137023 109059 137051
rect 109087 137023 109121 137051
rect 109149 137023 109184 137051
rect 109024 136989 109184 137023
rect 109024 136961 109059 136989
rect 109087 136961 109121 136989
rect 109149 136961 109184 136989
rect 109024 136944 109184 136961
rect 124384 137175 124544 137192
rect 124384 137147 124419 137175
rect 124447 137147 124481 137175
rect 124509 137147 124544 137175
rect 124384 137113 124544 137147
rect 124384 137085 124419 137113
rect 124447 137085 124481 137113
rect 124509 137085 124544 137113
rect 124384 137051 124544 137085
rect 124384 137023 124419 137051
rect 124447 137023 124481 137051
rect 124509 137023 124544 137051
rect 124384 136989 124544 137023
rect 124384 136961 124419 136989
rect 124447 136961 124481 136989
rect 124509 136961 124544 136989
rect 124384 136944 124544 136961
rect 139744 137175 139904 137192
rect 139744 137147 139779 137175
rect 139807 137147 139841 137175
rect 139869 137147 139904 137175
rect 139744 137113 139904 137147
rect 139744 137085 139779 137113
rect 139807 137085 139841 137113
rect 139869 137085 139904 137113
rect 139744 137051 139904 137085
rect 139744 137023 139779 137051
rect 139807 137023 139841 137051
rect 139869 137023 139904 137051
rect 139744 136989 139904 137023
rect 139744 136961 139779 136989
rect 139807 136961 139841 136989
rect 139869 136961 139904 136989
rect 139744 136944 139904 136961
rect 155104 137175 155264 137192
rect 155104 137147 155139 137175
rect 155167 137147 155201 137175
rect 155229 137147 155264 137175
rect 155104 137113 155264 137147
rect 155104 137085 155139 137113
rect 155167 137085 155201 137113
rect 155229 137085 155264 137113
rect 155104 137051 155264 137085
rect 155104 137023 155139 137051
rect 155167 137023 155201 137051
rect 155229 137023 155264 137051
rect 155104 136989 155264 137023
rect 155104 136961 155139 136989
rect 155167 136961 155201 136989
rect 155229 136961 155264 136989
rect 155104 136944 155264 136961
rect 170464 137175 170624 137192
rect 170464 137147 170499 137175
rect 170527 137147 170561 137175
rect 170589 137147 170624 137175
rect 170464 137113 170624 137147
rect 170464 137085 170499 137113
rect 170527 137085 170561 137113
rect 170589 137085 170624 137113
rect 170464 137051 170624 137085
rect 170464 137023 170499 137051
rect 170527 137023 170561 137051
rect 170589 137023 170624 137051
rect 170464 136989 170624 137023
rect 170464 136961 170499 136989
rect 170527 136961 170561 136989
rect 170589 136961 170624 136989
rect 170464 136944 170624 136961
rect 185824 137175 185984 137192
rect 185824 137147 185859 137175
rect 185887 137147 185921 137175
rect 185949 137147 185984 137175
rect 185824 137113 185984 137147
rect 185824 137085 185859 137113
rect 185887 137085 185921 137113
rect 185949 137085 185984 137113
rect 185824 137051 185984 137085
rect 185824 137023 185859 137051
rect 185887 137023 185921 137051
rect 185949 137023 185984 137051
rect 185824 136989 185984 137023
rect 185824 136961 185859 136989
rect 185887 136961 185921 136989
rect 185949 136961 185984 136989
rect 185824 136944 185984 136961
rect 201184 137175 201344 137192
rect 201184 137147 201219 137175
rect 201247 137147 201281 137175
rect 201309 137147 201344 137175
rect 201184 137113 201344 137147
rect 201184 137085 201219 137113
rect 201247 137085 201281 137113
rect 201309 137085 201344 137113
rect 201184 137051 201344 137085
rect 201184 137023 201219 137051
rect 201247 137023 201281 137051
rect 201309 137023 201344 137051
rect 201184 136989 201344 137023
rect 201184 136961 201219 136989
rect 201247 136961 201281 136989
rect 201309 136961 201344 136989
rect 201184 136944 201344 136961
rect 96729 131147 96777 131175
rect 96805 131147 96839 131175
rect 96867 131147 96901 131175
rect 96929 131147 96963 131175
rect 96991 131147 97039 131175
rect 96729 131113 97039 131147
rect 96729 131085 96777 131113
rect 96805 131085 96839 131113
rect 96867 131085 96901 131113
rect 96929 131085 96963 131113
rect 96991 131085 97039 131113
rect 96729 131051 97039 131085
rect 96729 131023 96777 131051
rect 96805 131023 96839 131051
rect 96867 131023 96901 131051
rect 96929 131023 96963 131051
rect 96991 131023 97039 131051
rect 204249 131175 204559 139961
rect 208864 140175 209024 140192
rect 208864 140147 208899 140175
rect 208927 140147 208961 140175
rect 208989 140147 209024 140175
rect 208864 140113 209024 140147
rect 208864 140085 208899 140113
rect 208927 140085 208961 140113
rect 208989 140085 209024 140113
rect 208864 140051 209024 140085
rect 208864 140023 208899 140051
rect 208927 140023 208961 140051
rect 208989 140023 209024 140051
rect 208864 139989 209024 140023
rect 208864 139961 208899 139989
rect 208927 139961 208961 139989
rect 208989 139961 209024 139989
rect 208864 139944 209024 139961
rect 216544 137175 216704 137192
rect 216544 137147 216579 137175
rect 216607 137147 216641 137175
rect 216669 137147 216704 137175
rect 216544 137113 216704 137147
rect 216544 137085 216579 137113
rect 216607 137085 216641 137113
rect 216669 137085 216704 137113
rect 216544 137051 216704 137085
rect 216544 137023 216579 137051
rect 216607 137023 216641 137051
rect 216669 137023 216704 137051
rect 216544 136989 216704 137023
rect 216544 136961 216579 136989
rect 216607 136961 216641 136989
rect 216669 136961 216704 136989
rect 216544 136944 216704 136961
rect 217749 137175 218059 145961
rect 217749 137147 217797 137175
rect 217825 137147 217859 137175
rect 217887 137147 217921 137175
rect 217949 137147 217983 137175
rect 218011 137147 218059 137175
rect 217749 137113 218059 137147
rect 217749 137085 217797 137113
rect 217825 137085 217859 137113
rect 217887 137085 217921 137113
rect 217949 137085 217983 137113
rect 218011 137085 218059 137113
rect 217749 137051 218059 137085
rect 217749 137023 217797 137051
rect 217825 137023 217859 137051
rect 217887 137023 217921 137051
rect 217949 137023 217983 137051
rect 218011 137023 218059 137051
rect 217749 136989 218059 137023
rect 217749 136961 217797 136989
rect 217825 136961 217859 136989
rect 217887 136961 217921 136989
rect 217949 136961 217983 136989
rect 218011 136961 218059 136989
rect 204249 131147 204297 131175
rect 204325 131147 204359 131175
rect 204387 131147 204421 131175
rect 204449 131147 204483 131175
rect 204511 131147 204559 131175
rect 204249 131113 204559 131147
rect 204249 131085 204297 131113
rect 204325 131085 204359 131113
rect 204387 131085 204421 131113
rect 204449 131085 204483 131113
rect 204511 131085 204559 131113
rect 204249 131051 204559 131085
rect 96729 130989 97039 131023
rect 96729 130961 96777 130989
rect 96805 130961 96839 130989
rect 96867 130961 96901 130989
rect 96929 130961 96963 130989
rect 96991 130961 97039 130989
rect 96729 122175 97039 130961
rect 112089 131014 112399 131025
rect 112089 130986 112137 131014
rect 112165 130986 112199 131014
rect 112227 130986 112261 131014
rect 112289 130986 112323 131014
rect 112351 130986 112399 131014
rect 112089 130952 112399 130986
rect 112089 130924 112137 130952
rect 112165 130924 112199 130952
rect 112227 130924 112261 130952
rect 112289 130924 112323 130952
rect 112351 130924 112399 130952
rect 107086 126714 107114 126719
rect 107086 126378 107114 126686
rect 107086 126345 107114 126350
rect 96729 122147 96777 122175
rect 96805 122147 96839 122175
rect 96867 122147 96901 122175
rect 96929 122147 96963 122175
rect 96991 122147 97039 122175
rect 96729 122113 97039 122147
rect 96729 122085 96777 122113
rect 96805 122085 96839 122113
rect 96867 122085 96901 122113
rect 96929 122085 96963 122113
rect 96991 122085 97039 122113
rect 96729 122051 97039 122085
rect 96729 122023 96777 122051
rect 96805 122023 96839 122051
rect 96867 122023 96901 122051
rect 96929 122023 96963 122051
rect 96991 122023 97039 122051
rect 96729 121989 97039 122023
rect 96729 121961 96777 121989
rect 96805 121961 96839 121989
rect 96867 121961 96901 121989
rect 96929 121961 96963 121989
rect 96991 121961 97039 121989
rect 96729 113175 97039 121961
rect 109904 122175 110064 122192
rect 109904 122147 109939 122175
rect 109967 122147 110001 122175
rect 110029 122147 110064 122175
rect 109904 122113 110064 122147
rect 109904 122085 109939 122113
rect 109967 122085 110001 122113
rect 110029 122085 110064 122113
rect 109904 122051 110064 122085
rect 109904 122023 109939 122051
rect 109967 122023 110001 122051
rect 110029 122023 110064 122051
rect 109904 121989 110064 122023
rect 109904 121961 109939 121989
rect 109967 121961 110001 121989
rect 110029 121961 110064 121989
rect 109904 121944 110064 121961
rect 112089 122175 112399 130924
rect 125589 128175 125899 131025
rect 125589 128147 125637 128175
rect 125665 128147 125699 128175
rect 125727 128147 125761 128175
rect 125789 128147 125823 128175
rect 125851 128147 125899 128175
rect 125589 128113 125899 128147
rect 125589 128085 125637 128113
rect 125665 128085 125699 128113
rect 125727 128085 125761 128113
rect 125789 128085 125823 128113
rect 125851 128085 125899 128113
rect 125589 128051 125899 128085
rect 125589 128023 125637 128051
rect 125665 128023 125699 128051
rect 125727 128023 125761 128051
rect 125789 128023 125823 128051
rect 125851 128023 125899 128051
rect 125589 127989 125899 128023
rect 125589 127961 125637 127989
rect 125665 127961 125699 127989
rect 125727 127961 125761 127989
rect 125789 127961 125823 127989
rect 125851 127961 125899 127989
rect 112089 122147 112137 122175
rect 112165 122147 112199 122175
rect 112227 122147 112261 122175
rect 112289 122147 112323 122175
rect 112351 122147 112399 122175
rect 112089 122113 112399 122147
rect 112089 122085 112137 122113
rect 112165 122085 112199 122113
rect 112227 122085 112261 122113
rect 112289 122085 112323 122113
rect 112351 122085 112399 122113
rect 112089 122051 112399 122085
rect 112089 122023 112137 122051
rect 112165 122023 112199 122051
rect 112227 122023 112261 122051
rect 112289 122023 112323 122051
rect 112351 122023 112399 122051
rect 112089 121989 112399 122023
rect 112089 121961 112137 121989
rect 112165 121961 112199 121989
rect 112227 121961 112261 121989
rect 112289 121961 112323 121989
rect 112351 121961 112399 121989
rect 112089 121415 112399 121961
rect 125264 122175 125424 122192
rect 125264 122147 125299 122175
rect 125327 122147 125361 122175
rect 125389 122147 125424 122175
rect 125264 122113 125424 122147
rect 125264 122085 125299 122113
rect 125327 122085 125361 122113
rect 125389 122085 125424 122113
rect 125264 122051 125424 122085
rect 125264 122023 125299 122051
rect 125327 122023 125361 122051
rect 125389 122023 125424 122051
rect 125264 121989 125424 122023
rect 125264 121961 125299 121989
rect 125327 121961 125361 121989
rect 125389 121961 125424 121989
rect 125264 121944 125424 121961
rect 102224 119175 102384 119192
rect 102224 119147 102259 119175
rect 102287 119147 102321 119175
rect 102349 119147 102384 119175
rect 102224 119113 102384 119147
rect 102224 119085 102259 119113
rect 102287 119085 102321 119113
rect 102349 119085 102384 119113
rect 102224 119051 102384 119085
rect 102224 119023 102259 119051
rect 102287 119023 102321 119051
rect 102349 119023 102384 119051
rect 102224 118989 102384 119023
rect 102224 118961 102259 118989
rect 102287 118961 102321 118989
rect 102349 118961 102384 118989
rect 102224 118944 102384 118961
rect 117584 119175 117744 119192
rect 117584 119147 117619 119175
rect 117647 119147 117681 119175
rect 117709 119147 117744 119175
rect 117584 119113 117744 119147
rect 117584 119085 117619 119113
rect 117647 119085 117681 119113
rect 117709 119085 117744 119113
rect 117584 119051 117744 119085
rect 117584 119023 117619 119051
rect 117647 119023 117681 119051
rect 117709 119023 117744 119051
rect 117584 118989 117744 119023
rect 117584 118961 117619 118989
rect 117647 118961 117681 118989
rect 117709 118961 117744 118989
rect 117584 118944 117744 118961
rect 125589 119175 125899 127961
rect 125589 119147 125637 119175
rect 125665 119147 125699 119175
rect 125727 119147 125761 119175
rect 125789 119147 125823 119175
rect 125851 119147 125899 119175
rect 125589 119113 125899 119147
rect 125589 119085 125637 119113
rect 125665 119085 125699 119113
rect 125727 119085 125761 119113
rect 125789 119085 125823 119113
rect 125851 119085 125899 119113
rect 125589 119051 125899 119085
rect 125589 119023 125637 119051
rect 125665 119023 125699 119051
rect 125727 119023 125761 119051
rect 125789 119023 125823 119051
rect 125851 119023 125899 119051
rect 125589 118989 125899 119023
rect 125589 118961 125637 118989
rect 125665 118961 125699 118989
rect 125727 118961 125761 118989
rect 125789 118961 125823 118989
rect 125851 118961 125899 118989
rect 96729 113147 96777 113175
rect 96805 113147 96839 113175
rect 96867 113147 96901 113175
rect 96929 113147 96963 113175
rect 96991 113147 97039 113175
rect 96729 113113 97039 113147
rect 96729 113085 96777 113113
rect 96805 113085 96839 113113
rect 96867 113085 96901 113113
rect 96929 113085 96963 113113
rect 96991 113085 97039 113113
rect 96729 113051 97039 113085
rect 96729 113023 96777 113051
rect 96805 113023 96839 113051
rect 96867 113023 96901 113051
rect 96929 113023 96963 113051
rect 96991 113023 97039 113051
rect 96729 112989 97039 113023
rect 96729 112961 96777 112989
rect 96805 112961 96839 112989
rect 96867 112961 96901 112989
rect 96929 112961 96963 112989
rect 96991 112961 97039 112989
rect 96729 104175 97039 112961
rect 109904 113175 110064 113192
rect 109904 113147 109939 113175
rect 109967 113147 110001 113175
rect 110029 113147 110064 113175
rect 109904 113113 110064 113147
rect 109904 113085 109939 113113
rect 109967 113085 110001 113113
rect 110029 113085 110064 113113
rect 109904 113051 110064 113085
rect 109904 113023 109939 113051
rect 109967 113023 110001 113051
rect 110029 113023 110064 113051
rect 109904 112989 110064 113023
rect 109904 112961 109939 112989
rect 109967 112961 110001 112989
rect 110029 112961 110064 112989
rect 109904 112944 110064 112961
rect 125264 113175 125424 113192
rect 125264 113147 125299 113175
rect 125327 113147 125361 113175
rect 125389 113147 125424 113175
rect 125264 113113 125424 113147
rect 125264 113085 125299 113113
rect 125327 113085 125361 113113
rect 125389 113085 125424 113113
rect 125264 113051 125424 113085
rect 125264 113023 125299 113051
rect 125327 113023 125361 113051
rect 125389 113023 125424 113051
rect 125264 112989 125424 113023
rect 125264 112961 125299 112989
rect 125327 112961 125361 112989
rect 125389 112961 125424 112989
rect 125264 112944 125424 112961
rect 102224 110175 102384 110192
rect 102224 110147 102259 110175
rect 102287 110147 102321 110175
rect 102349 110147 102384 110175
rect 102224 110113 102384 110147
rect 102224 110085 102259 110113
rect 102287 110085 102321 110113
rect 102349 110085 102384 110113
rect 102224 110051 102384 110085
rect 102224 110023 102259 110051
rect 102287 110023 102321 110051
rect 102349 110023 102384 110051
rect 102224 109989 102384 110023
rect 102224 109961 102259 109989
rect 102287 109961 102321 109989
rect 102349 109961 102384 109989
rect 102224 109944 102384 109961
rect 117584 110175 117744 110192
rect 117584 110147 117619 110175
rect 117647 110147 117681 110175
rect 117709 110147 117744 110175
rect 117584 110113 117744 110147
rect 117584 110085 117619 110113
rect 117647 110085 117681 110113
rect 117709 110085 117744 110113
rect 117584 110051 117744 110085
rect 117584 110023 117619 110051
rect 117647 110023 117681 110051
rect 117709 110023 117744 110051
rect 117584 109989 117744 110023
rect 117584 109961 117619 109989
rect 117647 109961 117681 109989
rect 117709 109961 117744 109989
rect 117584 109944 117744 109961
rect 125589 110175 125899 118961
rect 125589 110147 125637 110175
rect 125665 110147 125699 110175
rect 125727 110147 125761 110175
rect 125789 110147 125823 110175
rect 125851 110147 125899 110175
rect 125589 110113 125899 110147
rect 125589 110085 125637 110113
rect 125665 110085 125699 110113
rect 125727 110085 125761 110113
rect 125789 110085 125823 110113
rect 125851 110085 125899 110113
rect 125589 110051 125899 110085
rect 125589 110023 125637 110051
rect 125665 110023 125699 110051
rect 125727 110023 125761 110051
rect 125789 110023 125823 110051
rect 125851 110023 125899 110051
rect 125589 109989 125899 110023
rect 125589 109961 125637 109989
rect 125665 109961 125699 109989
rect 125727 109961 125761 109989
rect 125789 109961 125823 109989
rect 125851 109961 125899 109989
rect 96729 104147 96777 104175
rect 96805 104147 96839 104175
rect 96867 104147 96901 104175
rect 96929 104147 96963 104175
rect 96991 104147 97039 104175
rect 96729 104113 97039 104147
rect 96729 104085 96777 104113
rect 96805 104085 96839 104113
rect 96867 104085 96901 104113
rect 96929 104085 96963 104113
rect 96991 104085 97039 104113
rect 96729 104051 97039 104085
rect 96729 104023 96777 104051
rect 96805 104023 96839 104051
rect 96867 104023 96901 104051
rect 96929 104023 96963 104051
rect 96991 104023 97039 104051
rect 96729 103989 97039 104023
rect 96729 103961 96777 103989
rect 96805 103961 96839 103989
rect 96867 103961 96901 103989
rect 96929 103961 96963 103989
rect 96991 103961 97039 103989
rect 96729 95175 97039 103961
rect 109904 104175 110064 104192
rect 109904 104147 109939 104175
rect 109967 104147 110001 104175
rect 110029 104147 110064 104175
rect 109904 104113 110064 104147
rect 109904 104085 109939 104113
rect 109967 104085 110001 104113
rect 110029 104085 110064 104113
rect 109904 104051 110064 104085
rect 109904 104023 109939 104051
rect 109967 104023 110001 104051
rect 110029 104023 110064 104051
rect 109904 103989 110064 104023
rect 109904 103961 109939 103989
rect 109967 103961 110001 103989
rect 110029 103961 110064 103989
rect 109904 103944 110064 103961
rect 125264 104175 125424 104192
rect 125264 104147 125299 104175
rect 125327 104147 125361 104175
rect 125389 104147 125424 104175
rect 125264 104113 125424 104147
rect 125264 104085 125299 104113
rect 125327 104085 125361 104113
rect 125389 104085 125424 104113
rect 125264 104051 125424 104085
rect 125264 104023 125299 104051
rect 125327 104023 125361 104051
rect 125389 104023 125424 104051
rect 125264 103989 125424 104023
rect 125264 103961 125299 103989
rect 125327 103961 125361 103989
rect 125389 103961 125424 103989
rect 125264 103944 125424 103961
rect 102224 101175 102384 101192
rect 102224 101147 102259 101175
rect 102287 101147 102321 101175
rect 102349 101147 102384 101175
rect 102224 101113 102384 101147
rect 102224 101085 102259 101113
rect 102287 101085 102321 101113
rect 102349 101085 102384 101113
rect 102224 101051 102384 101085
rect 102224 101023 102259 101051
rect 102287 101023 102321 101051
rect 102349 101023 102384 101051
rect 102224 100989 102384 101023
rect 102224 100961 102259 100989
rect 102287 100961 102321 100989
rect 102349 100961 102384 100989
rect 102224 100944 102384 100961
rect 117584 101175 117744 101192
rect 117584 101147 117619 101175
rect 117647 101147 117681 101175
rect 117709 101147 117744 101175
rect 117584 101113 117744 101147
rect 117584 101085 117619 101113
rect 117647 101085 117681 101113
rect 117709 101085 117744 101113
rect 117584 101051 117744 101085
rect 117584 101023 117619 101051
rect 117647 101023 117681 101051
rect 117709 101023 117744 101051
rect 117584 100989 117744 101023
rect 117584 100961 117619 100989
rect 117647 100961 117681 100989
rect 117709 100961 117744 100989
rect 117584 100944 117744 100961
rect 125589 101175 125899 109961
rect 125589 101147 125637 101175
rect 125665 101147 125699 101175
rect 125727 101147 125761 101175
rect 125789 101147 125823 101175
rect 125851 101147 125899 101175
rect 125589 101113 125899 101147
rect 125589 101085 125637 101113
rect 125665 101085 125699 101113
rect 125727 101085 125761 101113
rect 125789 101085 125823 101113
rect 125851 101085 125899 101113
rect 125589 101051 125899 101085
rect 125589 101023 125637 101051
rect 125665 101023 125699 101051
rect 125727 101023 125761 101051
rect 125789 101023 125823 101051
rect 125851 101023 125899 101051
rect 125589 100989 125899 101023
rect 125589 100961 125637 100989
rect 125665 100961 125699 100989
rect 125727 100961 125761 100989
rect 125789 100961 125823 100989
rect 125851 100961 125899 100989
rect 96729 95147 96777 95175
rect 96805 95147 96839 95175
rect 96867 95147 96901 95175
rect 96929 95147 96963 95175
rect 96991 95147 97039 95175
rect 96729 95113 97039 95147
rect 96729 95085 96777 95113
rect 96805 95085 96839 95113
rect 96867 95085 96901 95113
rect 96929 95085 96963 95113
rect 96991 95085 97039 95113
rect 96729 95051 97039 95085
rect 96729 95023 96777 95051
rect 96805 95023 96839 95051
rect 96867 95023 96901 95051
rect 96929 95023 96963 95051
rect 96991 95023 97039 95051
rect 96729 94989 97039 95023
rect 96729 94961 96777 94989
rect 96805 94961 96839 94989
rect 96867 94961 96901 94989
rect 96929 94961 96963 94989
rect 96991 94961 97039 94989
rect 96729 86175 97039 94961
rect 96729 86147 96777 86175
rect 96805 86147 96839 86175
rect 96867 86147 96901 86175
rect 96929 86147 96963 86175
rect 96991 86147 97039 86175
rect 96729 86113 97039 86147
rect 96729 86085 96777 86113
rect 96805 86085 96839 86113
rect 96867 86085 96901 86113
rect 96929 86085 96963 86113
rect 96991 86085 97039 86113
rect 96729 86051 97039 86085
rect 96729 86023 96777 86051
rect 96805 86023 96839 86051
rect 96867 86023 96901 86051
rect 96929 86023 96963 86051
rect 96991 86023 97039 86051
rect 96729 85989 97039 86023
rect 96729 85961 96777 85989
rect 96805 85961 96839 85989
rect 96867 85961 96901 85989
rect 96929 85961 96963 85989
rect 96991 85961 97039 85989
rect 96729 77175 97039 85961
rect 96729 77147 96777 77175
rect 96805 77147 96839 77175
rect 96867 77147 96901 77175
rect 96929 77147 96963 77175
rect 96991 77147 97039 77175
rect 96729 77113 97039 77147
rect 96729 77085 96777 77113
rect 96805 77085 96839 77113
rect 96867 77085 96901 77113
rect 96929 77085 96963 77113
rect 96991 77085 97039 77113
rect 96729 77051 97039 77085
rect 96729 77023 96777 77051
rect 96805 77023 96839 77051
rect 96867 77023 96901 77051
rect 96929 77023 96963 77051
rect 96991 77023 97039 77051
rect 96729 76989 97039 77023
rect 96729 76961 96777 76989
rect 96805 76961 96839 76989
rect 96867 76961 96901 76989
rect 96929 76961 96963 76989
rect 96991 76961 97039 76989
rect 96729 68175 97039 76961
rect 96729 68147 96777 68175
rect 96805 68147 96839 68175
rect 96867 68147 96901 68175
rect 96929 68147 96963 68175
rect 96991 68147 97039 68175
rect 96729 68113 97039 68147
rect 96729 68085 96777 68113
rect 96805 68085 96839 68113
rect 96867 68085 96901 68113
rect 96929 68085 96963 68113
rect 96991 68085 97039 68113
rect 96729 68051 97039 68085
rect 96729 68023 96777 68051
rect 96805 68023 96839 68051
rect 96867 68023 96901 68051
rect 96929 68023 96963 68051
rect 96991 68023 97039 68051
rect 96729 67989 97039 68023
rect 96729 67961 96777 67989
rect 96805 67961 96839 67989
rect 96867 67961 96901 67989
rect 96929 67961 96963 67989
rect 96991 67961 97039 67989
rect 96729 59175 97039 67961
rect 96729 59147 96777 59175
rect 96805 59147 96839 59175
rect 96867 59147 96901 59175
rect 96929 59147 96963 59175
rect 96991 59147 97039 59175
rect 96729 59113 97039 59147
rect 96729 59085 96777 59113
rect 96805 59085 96839 59113
rect 96867 59085 96901 59113
rect 96929 59085 96963 59113
rect 96991 59085 97039 59113
rect 96729 59051 97039 59085
rect 96729 59023 96777 59051
rect 96805 59023 96839 59051
rect 96867 59023 96901 59051
rect 96929 59023 96963 59051
rect 96991 59023 97039 59051
rect 96729 58989 97039 59023
rect 96729 58961 96777 58989
rect 96805 58961 96839 58989
rect 96867 58961 96901 58989
rect 96929 58961 96963 58989
rect 96991 58961 97039 58989
rect 96729 50175 97039 58961
rect 96729 50147 96777 50175
rect 96805 50147 96839 50175
rect 96867 50147 96901 50175
rect 96929 50147 96963 50175
rect 96991 50147 97039 50175
rect 96729 50113 97039 50147
rect 96729 50085 96777 50113
rect 96805 50085 96839 50113
rect 96867 50085 96901 50113
rect 96929 50085 96963 50113
rect 96991 50085 97039 50113
rect 96729 50051 97039 50085
rect 96729 50023 96777 50051
rect 96805 50023 96839 50051
rect 96867 50023 96901 50051
rect 96929 50023 96963 50051
rect 96991 50023 97039 50051
rect 96729 49989 97039 50023
rect 96729 49961 96777 49989
rect 96805 49961 96839 49989
rect 96867 49961 96901 49989
rect 96929 49961 96963 49989
rect 96991 49961 97039 49989
rect 96729 41175 97039 49961
rect 96729 41147 96777 41175
rect 96805 41147 96839 41175
rect 96867 41147 96901 41175
rect 96929 41147 96963 41175
rect 96991 41147 97039 41175
rect 96729 41113 97039 41147
rect 96729 41085 96777 41113
rect 96805 41085 96839 41113
rect 96867 41085 96901 41113
rect 96929 41085 96963 41113
rect 96991 41085 97039 41113
rect 96729 41051 97039 41085
rect 96729 41023 96777 41051
rect 96805 41023 96839 41051
rect 96867 41023 96901 41051
rect 96929 41023 96963 41051
rect 96991 41023 97039 41051
rect 96729 40989 97039 41023
rect 96729 40961 96777 40989
rect 96805 40961 96839 40989
rect 96867 40961 96901 40989
rect 96929 40961 96963 40989
rect 96991 40961 97039 40989
rect 96729 32175 97039 40961
rect 96729 32147 96777 32175
rect 96805 32147 96839 32175
rect 96867 32147 96901 32175
rect 96929 32147 96963 32175
rect 96991 32147 97039 32175
rect 96729 32113 97039 32147
rect 96729 32085 96777 32113
rect 96805 32085 96839 32113
rect 96867 32085 96901 32113
rect 96929 32085 96963 32113
rect 96991 32085 97039 32113
rect 96729 32051 97039 32085
rect 96729 32023 96777 32051
rect 96805 32023 96839 32051
rect 96867 32023 96901 32051
rect 96929 32023 96963 32051
rect 96991 32023 97039 32051
rect 96729 31989 97039 32023
rect 96729 31961 96777 31989
rect 96805 31961 96839 31989
rect 96867 31961 96901 31989
rect 96929 31961 96963 31989
rect 96991 31961 97039 31989
rect 96729 23175 97039 31961
rect 96729 23147 96777 23175
rect 96805 23147 96839 23175
rect 96867 23147 96901 23175
rect 96929 23147 96963 23175
rect 96991 23147 97039 23175
rect 96729 23113 97039 23147
rect 96729 23085 96777 23113
rect 96805 23085 96839 23113
rect 96867 23085 96901 23113
rect 96929 23085 96963 23113
rect 96991 23085 97039 23113
rect 96729 23051 97039 23085
rect 96729 23023 96777 23051
rect 96805 23023 96839 23051
rect 96867 23023 96901 23051
rect 96929 23023 96963 23051
rect 96991 23023 97039 23051
rect 96729 22989 97039 23023
rect 96729 22961 96777 22989
rect 96805 22961 96839 22989
rect 96867 22961 96901 22989
rect 96929 22961 96963 22989
rect 96991 22961 97039 22989
rect 96729 14175 97039 22961
rect 96729 14147 96777 14175
rect 96805 14147 96839 14175
rect 96867 14147 96901 14175
rect 96929 14147 96963 14175
rect 96991 14147 97039 14175
rect 96729 14113 97039 14147
rect 96729 14085 96777 14113
rect 96805 14085 96839 14113
rect 96867 14085 96901 14113
rect 96929 14085 96963 14113
rect 96991 14085 97039 14113
rect 96729 14051 97039 14085
rect 96729 14023 96777 14051
rect 96805 14023 96839 14051
rect 96867 14023 96901 14051
rect 96929 14023 96963 14051
rect 96991 14023 97039 14051
rect 96729 13989 97039 14023
rect 96729 13961 96777 13989
rect 96805 13961 96839 13989
rect 96867 13961 96901 13989
rect 96929 13961 96963 13989
rect 96991 13961 97039 13989
rect 96729 5175 97039 13961
rect 96729 5147 96777 5175
rect 96805 5147 96839 5175
rect 96867 5147 96901 5175
rect 96929 5147 96963 5175
rect 96991 5147 97039 5175
rect 96729 5113 97039 5147
rect 96729 5085 96777 5113
rect 96805 5085 96839 5113
rect 96867 5085 96901 5113
rect 96929 5085 96963 5113
rect 96991 5085 97039 5113
rect 96729 5051 97039 5085
rect 96729 5023 96777 5051
rect 96805 5023 96839 5051
rect 96867 5023 96901 5051
rect 96929 5023 96963 5051
rect 96991 5023 97039 5051
rect 96729 4989 97039 5023
rect 96729 4961 96777 4989
rect 96805 4961 96839 4989
rect 96867 4961 96901 4989
rect 96929 4961 96963 4989
rect 96991 4961 97039 4989
rect 96729 -560 97039 4961
rect 96729 -588 96777 -560
rect 96805 -588 96839 -560
rect 96867 -588 96901 -560
rect 96929 -588 96963 -560
rect 96991 -588 97039 -560
rect 96729 -622 97039 -588
rect 96729 -650 96777 -622
rect 96805 -650 96839 -622
rect 96867 -650 96901 -622
rect 96929 -650 96963 -622
rect 96991 -650 97039 -622
rect 96729 -684 97039 -650
rect 96729 -712 96777 -684
rect 96805 -712 96839 -684
rect 96867 -712 96901 -684
rect 96929 -712 96963 -684
rect 96991 -712 97039 -684
rect 96729 -746 97039 -712
rect 96729 -774 96777 -746
rect 96805 -774 96839 -746
rect 96867 -774 96901 -746
rect 96929 -774 96963 -746
rect 96991 -774 97039 -746
rect 96729 -822 97039 -774
rect 110229 92175 110539 97761
rect 110229 92147 110277 92175
rect 110305 92147 110339 92175
rect 110367 92147 110401 92175
rect 110429 92147 110463 92175
rect 110491 92147 110539 92175
rect 110229 92113 110539 92147
rect 110229 92085 110277 92113
rect 110305 92085 110339 92113
rect 110367 92085 110401 92113
rect 110429 92085 110463 92113
rect 110491 92085 110539 92113
rect 110229 92051 110539 92085
rect 110229 92023 110277 92051
rect 110305 92023 110339 92051
rect 110367 92023 110401 92051
rect 110429 92023 110463 92051
rect 110491 92023 110539 92051
rect 110229 91989 110539 92023
rect 110229 91961 110277 91989
rect 110305 91961 110339 91989
rect 110367 91961 110401 91989
rect 110429 91961 110463 91989
rect 110491 91961 110539 91989
rect 110229 83175 110539 91961
rect 110229 83147 110277 83175
rect 110305 83147 110339 83175
rect 110367 83147 110401 83175
rect 110429 83147 110463 83175
rect 110491 83147 110539 83175
rect 110229 83113 110539 83147
rect 110229 83085 110277 83113
rect 110305 83085 110339 83113
rect 110367 83085 110401 83113
rect 110429 83085 110463 83113
rect 110491 83085 110539 83113
rect 110229 83051 110539 83085
rect 110229 83023 110277 83051
rect 110305 83023 110339 83051
rect 110367 83023 110401 83051
rect 110429 83023 110463 83051
rect 110491 83023 110539 83051
rect 110229 82989 110539 83023
rect 110229 82961 110277 82989
rect 110305 82961 110339 82989
rect 110367 82961 110401 82989
rect 110429 82961 110463 82989
rect 110491 82961 110539 82989
rect 110229 74175 110539 82961
rect 110229 74147 110277 74175
rect 110305 74147 110339 74175
rect 110367 74147 110401 74175
rect 110429 74147 110463 74175
rect 110491 74147 110539 74175
rect 110229 74113 110539 74147
rect 110229 74085 110277 74113
rect 110305 74085 110339 74113
rect 110367 74085 110401 74113
rect 110429 74085 110463 74113
rect 110491 74085 110539 74113
rect 110229 74051 110539 74085
rect 110229 74023 110277 74051
rect 110305 74023 110339 74051
rect 110367 74023 110401 74051
rect 110429 74023 110463 74051
rect 110491 74023 110539 74051
rect 110229 73989 110539 74023
rect 110229 73961 110277 73989
rect 110305 73961 110339 73989
rect 110367 73961 110401 73989
rect 110429 73961 110463 73989
rect 110491 73961 110539 73989
rect 110229 65175 110539 73961
rect 110229 65147 110277 65175
rect 110305 65147 110339 65175
rect 110367 65147 110401 65175
rect 110429 65147 110463 65175
rect 110491 65147 110539 65175
rect 110229 65113 110539 65147
rect 110229 65085 110277 65113
rect 110305 65085 110339 65113
rect 110367 65085 110401 65113
rect 110429 65085 110463 65113
rect 110491 65085 110539 65113
rect 110229 65051 110539 65085
rect 110229 65023 110277 65051
rect 110305 65023 110339 65051
rect 110367 65023 110401 65051
rect 110429 65023 110463 65051
rect 110491 65023 110539 65051
rect 110229 64989 110539 65023
rect 110229 64961 110277 64989
rect 110305 64961 110339 64989
rect 110367 64961 110401 64989
rect 110429 64961 110463 64989
rect 110491 64961 110539 64989
rect 110229 56175 110539 64961
rect 110229 56147 110277 56175
rect 110305 56147 110339 56175
rect 110367 56147 110401 56175
rect 110429 56147 110463 56175
rect 110491 56147 110539 56175
rect 110229 56113 110539 56147
rect 110229 56085 110277 56113
rect 110305 56085 110339 56113
rect 110367 56085 110401 56113
rect 110429 56085 110463 56113
rect 110491 56085 110539 56113
rect 110229 56051 110539 56085
rect 110229 56023 110277 56051
rect 110305 56023 110339 56051
rect 110367 56023 110401 56051
rect 110429 56023 110463 56051
rect 110491 56023 110539 56051
rect 110229 55989 110539 56023
rect 110229 55961 110277 55989
rect 110305 55961 110339 55989
rect 110367 55961 110401 55989
rect 110429 55961 110463 55989
rect 110491 55961 110539 55989
rect 110229 47175 110539 55961
rect 110229 47147 110277 47175
rect 110305 47147 110339 47175
rect 110367 47147 110401 47175
rect 110429 47147 110463 47175
rect 110491 47147 110539 47175
rect 110229 47113 110539 47147
rect 110229 47085 110277 47113
rect 110305 47085 110339 47113
rect 110367 47085 110401 47113
rect 110429 47085 110463 47113
rect 110491 47085 110539 47113
rect 110229 47051 110539 47085
rect 110229 47023 110277 47051
rect 110305 47023 110339 47051
rect 110367 47023 110401 47051
rect 110429 47023 110463 47051
rect 110491 47023 110539 47051
rect 110229 46989 110539 47023
rect 110229 46961 110277 46989
rect 110305 46961 110339 46989
rect 110367 46961 110401 46989
rect 110429 46961 110463 46989
rect 110491 46961 110539 46989
rect 110229 38175 110539 46961
rect 110229 38147 110277 38175
rect 110305 38147 110339 38175
rect 110367 38147 110401 38175
rect 110429 38147 110463 38175
rect 110491 38147 110539 38175
rect 110229 38113 110539 38147
rect 110229 38085 110277 38113
rect 110305 38085 110339 38113
rect 110367 38085 110401 38113
rect 110429 38085 110463 38113
rect 110491 38085 110539 38113
rect 110229 38051 110539 38085
rect 110229 38023 110277 38051
rect 110305 38023 110339 38051
rect 110367 38023 110401 38051
rect 110429 38023 110463 38051
rect 110491 38023 110539 38051
rect 110229 37989 110539 38023
rect 110229 37961 110277 37989
rect 110305 37961 110339 37989
rect 110367 37961 110401 37989
rect 110429 37961 110463 37989
rect 110491 37961 110539 37989
rect 110229 29175 110539 37961
rect 110229 29147 110277 29175
rect 110305 29147 110339 29175
rect 110367 29147 110401 29175
rect 110429 29147 110463 29175
rect 110491 29147 110539 29175
rect 110229 29113 110539 29147
rect 110229 29085 110277 29113
rect 110305 29085 110339 29113
rect 110367 29085 110401 29113
rect 110429 29085 110463 29113
rect 110491 29085 110539 29113
rect 110229 29051 110539 29085
rect 110229 29023 110277 29051
rect 110305 29023 110339 29051
rect 110367 29023 110401 29051
rect 110429 29023 110463 29051
rect 110491 29023 110539 29051
rect 110229 28989 110539 29023
rect 110229 28961 110277 28989
rect 110305 28961 110339 28989
rect 110367 28961 110401 28989
rect 110429 28961 110463 28989
rect 110491 28961 110539 28989
rect 110229 20175 110539 28961
rect 110229 20147 110277 20175
rect 110305 20147 110339 20175
rect 110367 20147 110401 20175
rect 110429 20147 110463 20175
rect 110491 20147 110539 20175
rect 110229 20113 110539 20147
rect 110229 20085 110277 20113
rect 110305 20085 110339 20113
rect 110367 20085 110401 20113
rect 110429 20085 110463 20113
rect 110491 20085 110539 20113
rect 110229 20051 110539 20085
rect 110229 20023 110277 20051
rect 110305 20023 110339 20051
rect 110367 20023 110401 20051
rect 110429 20023 110463 20051
rect 110491 20023 110539 20051
rect 110229 19989 110539 20023
rect 110229 19961 110277 19989
rect 110305 19961 110339 19989
rect 110367 19961 110401 19989
rect 110429 19961 110463 19989
rect 110491 19961 110539 19989
rect 110229 11175 110539 19961
rect 110229 11147 110277 11175
rect 110305 11147 110339 11175
rect 110367 11147 110401 11175
rect 110429 11147 110463 11175
rect 110491 11147 110539 11175
rect 110229 11113 110539 11147
rect 110229 11085 110277 11113
rect 110305 11085 110339 11113
rect 110367 11085 110401 11113
rect 110429 11085 110463 11113
rect 110491 11085 110539 11113
rect 110229 11051 110539 11085
rect 110229 11023 110277 11051
rect 110305 11023 110339 11051
rect 110367 11023 110401 11051
rect 110429 11023 110463 11051
rect 110491 11023 110539 11051
rect 110229 10989 110539 11023
rect 110229 10961 110277 10989
rect 110305 10961 110339 10989
rect 110367 10961 110401 10989
rect 110429 10961 110463 10989
rect 110491 10961 110539 10989
rect 110229 2175 110539 10961
rect 110229 2147 110277 2175
rect 110305 2147 110339 2175
rect 110367 2147 110401 2175
rect 110429 2147 110463 2175
rect 110491 2147 110539 2175
rect 110229 2113 110539 2147
rect 110229 2085 110277 2113
rect 110305 2085 110339 2113
rect 110367 2085 110401 2113
rect 110429 2085 110463 2113
rect 110491 2085 110539 2113
rect 110229 2051 110539 2085
rect 110229 2023 110277 2051
rect 110305 2023 110339 2051
rect 110367 2023 110401 2051
rect 110429 2023 110463 2051
rect 110491 2023 110539 2051
rect 110229 1989 110539 2023
rect 110229 1961 110277 1989
rect 110305 1961 110339 1989
rect 110367 1961 110401 1989
rect 110429 1961 110463 1989
rect 110491 1961 110539 1989
rect 110229 -80 110539 1961
rect 110229 -108 110277 -80
rect 110305 -108 110339 -80
rect 110367 -108 110401 -80
rect 110429 -108 110463 -80
rect 110491 -108 110539 -80
rect 110229 -142 110539 -108
rect 110229 -170 110277 -142
rect 110305 -170 110339 -142
rect 110367 -170 110401 -142
rect 110429 -170 110463 -142
rect 110491 -170 110539 -142
rect 110229 -204 110539 -170
rect 110229 -232 110277 -204
rect 110305 -232 110339 -204
rect 110367 -232 110401 -204
rect 110429 -232 110463 -204
rect 110491 -232 110539 -204
rect 110229 -266 110539 -232
rect 110229 -294 110277 -266
rect 110305 -294 110339 -266
rect 110367 -294 110401 -266
rect 110429 -294 110463 -266
rect 110491 -294 110539 -266
rect 110229 -822 110539 -294
rect 112089 95175 112399 97761
rect 112089 95147 112137 95175
rect 112165 95147 112199 95175
rect 112227 95147 112261 95175
rect 112289 95147 112323 95175
rect 112351 95147 112399 95175
rect 112089 95113 112399 95147
rect 112089 95085 112137 95113
rect 112165 95085 112199 95113
rect 112227 95085 112261 95113
rect 112289 95085 112323 95113
rect 112351 95085 112399 95113
rect 112089 95051 112399 95085
rect 112089 95023 112137 95051
rect 112165 95023 112199 95051
rect 112227 95023 112261 95051
rect 112289 95023 112323 95051
rect 112351 95023 112399 95051
rect 112089 94989 112399 95023
rect 112089 94961 112137 94989
rect 112165 94961 112199 94989
rect 112227 94961 112261 94989
rect 112289 94961 112323 94989
rect 112351 94961 112399 94989
rect 112089 86175 112399 94961
rect 112089 86147 112137 86175
rect 112165 86147 112199 86175
rect 112227 86147 112261 86175
rect 112289 86147 112323 86175
rect 112351 86147 112399 86175
rect 112089 86113 112399 86147
rect 112089 86085 112137 86113
rect 112165 86085 112199 86113
rect 112227 86085 112261 86113
rect 112289 86085 112323 86113
rect 112351 86085 112399 86113
rect 112089 86051 112399 86085
rect 112089 86023 112137 86051
rect 112165 86023 112199 86051
rect 112227 86023 112261 86051
rect 112289 86023 112323 86051
rect 112351 86023 112399 86051
rect 112089 85989 112399 86023
rect 112089 85961 112137 85989
rect 112165 85961 112199 85989
rect 112227 85961 112261 85989
rect 112289 85961 112323 85989
rect 112351 85961 112399 85989
rect 112089 77175 112399 85961
rect 112089 77147 112137 77175
rect 112165 77147 112199 77175
rect 112227 77147 112261 77175
rect 112289 77147 112323 77175
rect 112351 77147 112399 77175
rect 112089 77113 112399 77147
rect 112089 77085 112137 77113
rect 112165 77085 112199 77113
rect 112227 77085 112261 77113
rect 112289 77085 112323 77113
rect 112351 77085 112399 77113
rect 112089 77051 112399 77085
rect 112089 77023 112137 77051
rect 112165 77023 112199 77051
rect 112227 77023 112261 77051
rect 112289 77023 112323 77051
rect 112351 77023 112399 77051
rect 112089 76989 112399 77023
rect 112089 76961 112137 76989
rect 112165 76961 112199 76989
rect 112227 76961 112261 76989
rect 112289 76961 112323 76989
rect 112351 76961 112399 76989
rect 112089 68175 112399 76961
rect 112089 68147 112137 68175
rect 112165 68147 112199 68175
rect 112227 68147 112261 68175
rect 112289 68147 112323 68175
rect 112351 68147 112399 68175
rect 112089 68113 112399 68147
rect 112089 68085 112137 68113
rect 112165 68085 112199 68113
rect 112227 68085 112261 68113
rect 112289 68085 112323 68113
rect 112351 68085 112399 68113
rect 112089 68051 112399 68085
rect 112089 68023 112137 68051
rect 112165 68023 112199 68051
rect 112227 68023 112261 68051
rect 112289 68023 112323 68051
rect 112351 68023 112399 68051
rect 112089 67989 112399 68023
rect 112089 67961 112137 67989
rect 112165 67961 112199 67989
rect 112227 67961 112261 67989
rect 112289 67961 112323 67989
rect 112351 67961 112399 67989
rect 112089 59175 112399 67961
rect 112089 59147 112137 59175
rect 112165 59147 112199 59175
rect 112227 59147 112261 59175
rect 112289 59147 112323 59175
rect 112351 59147 112399 59175
rect 112089 59113 112399 59147
rect 112089 59085 112137 59113
rect 112165 59085 112199 59113
rect 112227 59085 112261 59113
rect 112289 59085 112323 59113
rect 112351 59085 112399 59113
rect 112089 59051 112399 59085
rect 112089 59023 112137 59051
rect 112165 59023 112199 59051
rect 112227 59023 112261 59051
rect 112289 59023 112323 59051
rect 112351 59023 112399 59051
rect 112089 58989 112399 59023
rect 112089 58961 112137 58989
rect 112165 58961 112199 58989
rect 112227 58961 112261 58989
rect 112289 58961 112323 58989
rect 112351 58961 112399 58989
rect 112089 50175 112399 58961
rect 112089 50147 112137 50175
rect 112165 50147 112199 50175
rect 112227 50147 112261 50175
rect 112289 50147 112323 50175
rect 112351 50147 112399 50175
rect 112089 50113 112399 50147
rect 112089 50085 112137 50113
rect 112165 50085 112199 50113
rect 112227 50085 112261 50113
rect 112289 50085 112323 50113
rect 112351 50085 112399 50113
rect 112089 50051 112399 50085
rect 112089 50023 112137 50051
rect 112165 50023 112199 50051
rect 112227 50023 112261 50051
rect 112289 50023 112323 50051
rect 112351 50023 112399 50051
rect 112089 49989 112399 50023
rect 112089 49961 112137 49989
rect 112165 49961 112199 49989
rect 112227 49961 112261 49989
rect 112289 49961 112323 49989
rect 112351 49961 112399 49989
rect 112089 41175 112399 49961
rect 112089 41147 112137 41175
rect 112165 41147 112199 41175
rect 112227 41147 112261 41175
rect 112289 41147 112323 41175
rect 112351 41147 112399 41175
rect 112089 41113 112399 41147
rect 112089 41085 112137 41113
rect 112165 41085 112199 41113
rect 112227 41085 112261 41113
rect 112289 41085 112323 41113
rect 112351 41085 112399 41113
rect 112089 41051 112399 41085
rect 112089 41023 112137 41051
rect 112165 41023 112199 41051
rect 112227 41023 112261 41051
rect 112289 41023 112323 41051
rect 112351 41023 112399 41051
rect 112089 40989 112399 41023
rect 112089 40961 112137 40989
rect 112165 40961 112199 40989
rect 112227 40961 112261 40989
rect 112289 40961 112323 40989
rect 112351 40961 112399 40989
rect 112089 32175 112399 40961
rect 112089 32147 112137 32175
rect 112165 32147 112199 32175
rect 112227 32147 112261 32175
rect 112289 32147 112323 32175
rect 112351 32147 112399 32175
rect 112089 32113 112399 32147
rect 112089 32085 112137 32113
rect 112165 32085 112199 32113
rect 112227 32085 112261 32113
rect 112289 32085 112323 32113
rect 112351 32085 112399 32113
rect 112089 32051 112399 32085
rect 112089 32023 112137 32051
rect 112165 32023 112199 32051
rect 112227 32023 112261 32051
rect 112289 32023 112323 32051
rect 112351 32023 112399 32051
rect 112089 31989 112399 32023
rect 112089 31961 112137 31989
rect 112165 31961 112199 31989
rect 112227 31961 112261 31989
rect 112289 31961 112323 31989
rect 112351 31961 112399 31989
rect 112089 23175 112399 31961
rect 112089 23147 112137 23175
rect 112165 23147 112199 23175
rect 112227 23147 112261 23175
rect 112289 23147 112323 23175
rect 112351 23147 112399 23175
rect 112089 23113 112399 23147
rect 112089 23085 112137 23113
rect 112165 23085 112199 23113
rect 112227 23085 112261 23113
rect 112289 23085 112323 23113
rect 112351 23085 112399 23113
rect 112089 23051 112399 23085
rect 112089 23023 112137 23051
rect 112165 23023 112199 23051
rect 112227 23023 112261 23051
rect 112289 23023 112323 23051
rect 112351 23023 112399 23051
rect 112089 22989 112399 23023
rect 112089 22961 112137 22989
rect 112165 22961 112199 22989
rect 112227 22961 112261 22989
rect 112289 22961 112323 22989
rect 112351 22961 112399 22989
rect 112089 14175 112399 22961
rect 112089 14147 112137 14175
rect 112165 14147 112199 14175
rect 112227 14147 112261 14175
rect 112289 14147 112323 14175
rect 112351 14147 112399 14175
rect 112089 14113 112399 14147
rect 112089 14085 112137 14113
rect 112165 14085 112199 14113
rect 112227 14085 112261 14113
rect 112289 14085 112323 14113
rect 112351 14085 112399 14113
rect 112089 14051 112399 14085
rect 112089 14023 112137 14051
rect 112165 14023 112199 14051
rect 112227 14023 112261 14051
rect 112289 14023 112323 14051
rect 112351 14023 112399 14051
rect 112089 13989 112399 14023
rect 112089 13961 112137 13989
rect 112165 13961 112199 13989
rect 112227 13961 112261 13989
rect 112289 13961 112323 13989
rect 112351 13961 112399 13989
rect 112089 5175 112399 13961
rect 112089 5147 112137 5175
rect 112165 5147 112199 5175
rect 112227 5147 112261 5175
rect 112289 5147 112323 5175
rect 112351 5147 112399 5175
rect 112089 5113 112399 5147
rect 112089 5085 112137 5113
rect 112165 5085 112199 5113
rect 112227 5085 112261 5113
rect 112289 5085 112323 5113
rect 112351 5085 112399 5113
rect 112089 5051 112399 5085
rect 112089 5023 112137 5051
rect 112165 5023 112199 5051
rect 112227 5023 112261 5051
rect 112289 5023 112323 5051
rect 112351 5023 112399 5051
rect 112089 4989 112399 5023
rect 112089 4961 112137 4989
rect 112165 4961 112199 4989
rect 112227 4961 112261 4989
rect 112289 4961 112323 4989
rect 112351 4961 112399 4989
rect 112089 -560 112399 4961
rect 112089 -588 112137 -560
rect 112165 -588 112199 -560
rect 112227 -588 112261 -560
rect 112289 -588 112323 -560
rect 112351 -588 112399 -560
rect 112089 -622 112399 -588
rect 112089 -650 112137 -622
rect 112165 -650 112199 -622
rect 112227 -650 112261 -622
rect 112289 -650 112323 -622
rect 112351 -650 112399 -622
rect 112089 -684 112399 -650
rect 112089 -712 112137 -684
rect 112165 -712 112199 -684
rect 112227 -712 112261 -684
rect 112289 -712 112323 -684
rect 112351 -712 112399 -684
rect 112089 -746 112399 -712
rect 112089 -774 112137 -746
rect 112165 -774 112199 -746
rect 112227 -774 112261 -746
rect 112289 -774 112323 -746
rect 112351 -774 112399 -746
rect 112089 -822 112399 -774
rect 125589 92175 125899 100961
rect 125589 92147 125637 92175
rect 125665 92147 125699 92175
rect 125727 92147 125761 92175
rect 125789 92147 125823 92175
rect 125851 92147 125899 92175
rect 125589 92113 125899 92147
rect 125589 92085 125637 92113
rect 125665 92085 125699 92113
rect 125727 92085 125761 92113
rect 125789 92085 125823 92113
rect 125851 92085 125899 92113
rect 125589 92051 125899 92085
rect 125589 92023 125637 92051
rect 125665 92023 125699 92051
rect 125727 92023 125761 92051
rect 125789 92023 125823 92051
rect 125851 92023 125899 92051
rect 125589 91989 125899 92023
rect 125589 91961 125637 91989
rect 125665 91961 125699 91989
rect 125727 91961 125761 91989
rect 125789 91961 125823 91989
rect 125851 91961 125899 91989
rect 125589 83175 125899 91961
rect 125589 83147 125637 83175
rect 125665 83147 125699 83175
rect 125727 83147 125761 83175
rect 125789 83147 125823 83175
rect 125851 83147 125899 83175
rect 125589 83113 125899 83147
rect 125589 83085 125637 83113
rect 125665 83085 125699 83113
rect 125727 83085 125761 83113
rect 125789 83085 125823 83113
rect 125851 83085 125899 83113
rect 125589 83051 125899 83085
rect 125589 83023 125637 83051
rect 125665 83023 125699 83051
rect 125727 83023 125761 83051
rect 125789 83023 125823 83051
rect 125851 83023 125899 83051
rect 125589 82989 125899 83023
rect 125589 82961 125637 82989
rect 125665 82961 125699 82989
rect 125727 82961 125761 82989
rect 125789 82961 125823 82989
rect 125851 82961 125899 82989
rect 125589 74175 125899 82961
rect 125589 74147 125637 74175
rect 125665 74147 125699 74175
rect 125727 74147 125761 74175
rect 125789 74147 125823 74175
rect 125851 74147 125899 74175
rect 125589 74113 125899 74147
rect 125589 74085 125637 74113
rect 125665 74085 125699 74113
rect 125727 74085 125761 74113
rect 125789 74085 125823 74113
rect 125851 74085 125899 74113
rect 125589 74051 125899 74085
rect 125589 74023 125637 74051
rect 125665 74023 125699 74051
rect 125727 74023 125761 74051
rect 125789 74023 125823 74051
rect 125851 74023 125899 74051
rect 125589 73989 125899 74023
rect 125589 73961 125637 73989
rect 125665 73961 125699 73989
rect 125727 73961 125761 73989
rect 125789 73961 125823 73989
rect 125851 73961 125899 73989
rect 125589 65175 125899 73961
rect 125589 65147 125637 65175
rect 125665 65147 125699 65175
rect 125727 65147 125761 65175
rect 125789 65147 125823 65175
rect 125851 65147 125899 65175
rect 125589 65113 125899 65147
rect 125589 65085 125637 65113
rect 125665 65085 125699 65113
rect 125727 65085 125761 65113
rect 125789 65085 125823 65113
rect 125851 65085 125899 65113
rect 125589 65051 125899 65085
rect 125589 65023 125637 65051
rect 125665 65023 125699 65051
rect 125727 65023 125761 65051
rect 125789 65023 125823 65051
rect 125851 65023 125899 65051
rect 125589 64989 125899 65023
rect 125589 64961 125637 64989
rect 125665 64961 125699 64989
rect 125727 64961 125761 64989
rect 125789 64961 125823 64989
rect 125851 64961 125899 64989
rect 125589 56175 125899 64961
rect 125589 56147 125637 56175
rect 125665 56147 125699 56175
rect 125727 56147 125761 56175
rect 125789 56147 125823 56175
rect 125851 56147 125899 56175
rect 125589 56113 125899 56147
rect 125589 56085 125637 56113
rect 125665 56085 125699 56113
rect 125727 56085 125761 56113
rect 125789 56085 125823 56113
rect 125851 56085 125899 56113
rect 125589 56051 125899 56085
rect 125589 56023 125637 56051
rect 125665 56023 125699 56051
rect 125727 56023 125761 56051
rect 125789 56023 125823 56051
rect 125851 56023 125899 56051
rect 125589 55989 125899 56023
rect 125589 55961 125637 55989
rect 125665 55961 125699 55989
rect 125727 55961 125761 55989
rect 125789 55961 125823 55989
rect 125851 55961 125899 55989
rect 125589 47175 125899 55961
rect 125589 47147 125637 47175
rect 125665 47147 125699 47175
rect 125727 47147 125761 47175
rect 125789 47147 125823 47175
rect 125851 47147 125899 47175
rect 125589 47113 125899 47147
rect 125589 47085 125637 47113
rect 125665 47085 125699 47113
rect 125727 47085 125761 47113
rect 125789 47085 125823 47113
rect 125851 47085 125899 47113
rect 125589 47051 125899 47085
rect 125589 47023 125637 47051
rect 125665 47023 125699 47051
rect 125727 47023 125761 47051
rect 125789 47023 125823 47051
rect 125851 47023 125899 47051
rect 125589 46989 125899 47023
rect 125589 46961 125637 46989
rect 125665 46961 125699 46989
rect 125727 46961 125761 46989
rect 125789 46961 125823 46989
rect 125851 46961 125899 46989
rect 125589 38175 125899 46961
rect 125589 38147 125637 38175
rect 125665 38147 125699 38175
rect 125727 38147 125761 38175
rect 125789 38147 125823 38175
rect 125851 38147 125899 38175
rect 125589 38113 125899 38147
rect 125589 38085 125637 38113
rect 125665 38085 125699 38113
rect 125727 38085 125761 38113
rect 125789 38085 125823 38113
rect 125851 38085 125899 38113
rect 125589 38051 125899 38085
rect 125589 38023 125637 38051
rect 125665 38023 125699 38051
rect 125727 38023 125761 38051
rect 125789 38023 125823 38051
rect 125851 38023 125899 38051
rect 125589 37989 125899 38023
rect 125589 37961 125637 37989
rect 125665 37961 125699 37989
rect 125727 37961 125761 37989
rect 125789 37961 125823 37989
rect 125851 37961 125899 37989
rect 125589 29175 125899 37961
rect 125589 29147 125637 29175
rect 125665 29147 125699 29175
rect 125727 29147 125761 29175
rect 125789 29147 125823 29175
rect 125851 29147 125899 29175
rect 125589 29113 125899 29147
rect 125589 29085 125637 29113
rect 125665 29085 125699 29113
rect 125727 29085 125761 29113
rect 125789 29085 125823 29113
rect 125851 29085 125899 29113
rect 125589 29051 125899 29085
rect 125589 29023 125637 29051
rect 125665 29023 125699 29051
rect 125727 29023 125761 29051
rect 125789 29023 125823 29051
rect 125851 29023 125899 29051
rect 125589 28989 125899 29023
rect 125589 28961 125637 28989
rect 125665 28961 125699 28989
rect 125727 28961 125761 28989
rect 125789 28961 125823 28989
rect 125851 28961 125899 28989
rect 125589 20175 125899 28961
rect 125589 20147 125637 20175
rect 125665 20147 125699 20175
rect 125727 20147 125761 20175
rect 125789 20147 125823 20175
rect 125851 20147 125899 20175
rect 125589 20113 125899 20147
rect 125589 20085 125637 20113
rect 125665 20085 125699 20113
rect 125727 20085 125761 20113
rect 125789 20085 125823 20113
rect 125851 20085 125899 20113
rect 125589 20051 125899 20085
rect 125589 20023 125637 20051
rect 125665 20023 125699 20051
rect 125727 20023 125761 20051
rect 125789 20023 125823 20051
rect 125851 20023 125899 20051
rect 125589 19989 125899 20023
rect 125589 19961 125637 19989
rect 125665 19961 125699 19989
rect 125727 19961 125761 19989
rect 125789 19961 125823 19989
rect 125851 19961 125899 19989
rect 125589 11175 125899 19961
rect 125589 11147 125637 11175
rect 125665 11147 125699 11175
rect 125727 11147 125761 11175
rect 125789 11147 125823 11175
rect 125851 11147 125899 11175
rect 125589 11113 125899 11147
rect 125589 11085 125637 11113
rect 125665 11085 125699 11113
rect 125727 11085 125761 11113
rect 125789 11085 125823 11113
rect 125851 11085 125899 11113
rect 125589 11051 125899 11085
rect 125589 11023 125637 11051
rect 125665 11023 125699 11051
rect 125727 11023 125761 11051
rect 125789 11023 125823 11051
rect 125851 11023 125899 11051
rect 125589 10989 125899 11023
rect 125589 10961 125637 10989
rect 125665 10961 125699 10989
rect 125727 10961 125761 10989
rect 125789 10961 125823 10989
rect 125851 10961 125899 10989
rect 125589 2175 125899 10961
rect 125589 2147 125637 2175
rect 125665 2147 125699 2175
rect 125727 2147 125761 2175
rect 125789 2147 125823 2175
rect 125851 2147 125899 2175
rect 125589 2113 125899 2147
rect 125589 2085 125637 2113
rect 125665 2085 125699 2113
rect 125727 2085 125761 2113
rect 125789 2085 125823 2113
rect 125851 2085 125899 2113
rect 125589 2051 125899 2085
rect 125589 2023 125637 2051
rect 125665 2023 125699 2051
rect 125727 2023 125761 2051
rect 125789 2023 125823 2051
rect 125851 2023 125899 2051
rect 125589 1989 125899 2023
rect 125589 1961 125637 1989
rect 125665 1961 125699 1989
rect 125727 1961 125761 1989
rect 125789 1961 125823 1989
rect 125851 1961 125899 1989
rect 125589 -80 125899 1961
rect 125589 -108 125637 -80
rect 125665 -108 125699 -80
rect 125727 -108 125761 -80
rect 125789 -108 125823 -80
rect 125851 -108 125899 -80
rect 125589 -142 125899 -108
rect 125589 -170 125637 -142
rect 125665 -170 125699 -142
rect 125727 -170 125761 -142
rect 125789 -170 125823 -142
rect 125851 -170 125899 -142
rect 125589 -204 125899 -170
rect 125589 -232 125637 -204
rect 125665 -232 125699 -204
rect 125727 -232 125761 -204
rect 125789 -232 125823 -204
rect 125851 -232 125899 -204
rect 125589 -266 125899 -232
rect 125589 -294 125637 -266
rect 125665 -294 125699 -266
rect 125727 -294 125761 -266
rect 125789 -294 125823 -266
rect 125851 -294 125899 -266
rect 125589 -822 125899 -294
rect 127449 131014 127759 131025
rect 127449 130986 127497 131014
rect 127525 130986 127559 131014
rect 127587 130986 127621 131014
rect 127649 130986 127683 131014
rect 127711 130986 127759 131014
rect 127449 130952 127759 130986
rect 127449 130924 127497 130952
rect 127525 130924 127559 130952
rect 127587 130924 127621 130952
rect 127649 130924 127683 130952
rect 127711 130924 127759 130952
rect 127449 122175 127759 130924
rect 127449 122147 127497 122175
rect 127525 122147 127559 122175
rect 127587 122147 127621 122175
rect 127649 122147 127683 122175
rect 127711 122147 127759 122175
rect 127449 122113 127759 122147
rect 127449 122085 127497 122113
rect 127525 122085 127559 122113
rect 127587 122085 127621 122113
rect 127649 122085 127683 122113
rect 127711 122085 127759 122113
rect 127449 122051 127759 122085
rect 127449 122023 127497 122051
rect 127525 122023 127559 122051
rect 127587 122023 127621 122051
rect 127649 122023 127683 122051
rect 127711 122023 127759 122051
rect 127449 121989 127759 122023
rect 127449 121961 127497 121989
rect 127525 121961 127559 121989
rect 127587 121961 127621 121989
rect 127649 121961 127683 121989
rect 127711 121961 127759 121989
rect 127449 113175 127759 121961
rect 127449 113147 127497 113175
rect 127525 113147 127559 113175
rect 127587 113147 127621 113175
rect 127649 113147 127683 113175
rect 127711 113147 127759 113175
rect 127449 113113 127759 113147
rect 127449 113085 127497 113113
rect 127525 113085 127559 113113
rect 127587 113085 127621 113113
rect 127649 113085 127683 113113
rect 127711 113085 127759 113113
rect 127449 113051 127759 113085
rect 127449 113023 127497 113051
rect 127525 113023 127559 113051
rect 127587 113023 127621 113051
rect 127649 113023 127683 113051
rect 127711 113023 127759 113051
rect 127449 112989 127759 113023
rect 127449 112961 127497 112989
rect 127525 112961 127559 112989
rect 127587 112961 127621 112989
rect 127649 112961 127683 112989
rect 127711 112961 127759 112989
rect 127449 104175 127759 112961
rect 127449 104147 127497 104175
rect 127525 104147 127559 104175
rect 127587 104147 127621 104175
rect 127649 104147 127683 104175
rect 127711 104147 127759 104175
rect 127449 104113 127759 104147
rect 127449 104085 127497 104113
rect 127525 104085 127559 104113
rect 127587 104085 127621 104113
rect 127649 104085 127683 104113
rect 127711 104085 127759 104113
rect 127449 104051 127759 104085
rect 127449 104023 127497 104051
rect 127525 104023 127559 104051
rect 127587 104023 127621 104051
rect 127649 104023 127683 104051
rect 127711 104023 127759 104051
rect 127449 103989 127759 104023
rect 127449 103961 127497 103989
rect 127525 103961 127559 103989
rect 127587 103961 127621 103989
rect 127649 103961 127683 103989
rect 127711 103961 127759 103989
rect 127449 95175 127759 103961
rect 127449 95147 127497 95175
rect 127525 95147 127559 95175
rect 127587 95147 127621 95175
rect 127649 95147 127683 95175
rect 127711 95147 127759 95175
rect 127449 95113 127759 95147
rect 127449 95085 127497 95113
rect 127525 95085 127559 95113
rect 127587 95085 127621 95113
rect 127649 95085 127683 95113
rect 127711 95085 127759 95113
rect 127449 95051 127759 95085
rect 127449 95023 127497 95051
rect 127525 95023 127559 95051
rect 127587 95023 127621 95051
rect 127649 95023 127683 95051
rect 127711 95023 127759 95051
rect 127449 94989 127759 95023
rect 127449 94961 127497 94989
rect 127525 94961 127559 94989
rect 127587 94961 127621 94989
rect 127649 94961 127683 94989
rect 127711 94961 127759 94989
rect 127449 86175 127759 94961
rect 127449 86147 127497 86175
rect 127525 86147 127559 86175
rect 127587 86147 127621 86175
rect 127649 86147 127683 86175
rect 127711 86147 127759 86175
rect 127449 86113 127759 86147
rect 127449 86085 127497 86113
rect 127525 86085 127559 86113
rect 127587 86085 127621 86113
rect 127649 86085 127683 86113
rect 127711 86085 127759 86113
rect 127449 86051 127759 86085
rect 127449 86023 127497 86051
rect 127525 86023 127559 86051
rect 127587 86023 127621 86051
rect 127649 86023 127683 86051
rect 127711 86023 127759 86051
rect 127449 85989 127759 86023
rect 127449 85961 127497 85989
rect 127525 85961 127559 85989
rect 127587 85961 127621 85989
rect 127649 85961 127683 85989
rect 127711 85961 127759 85989
rect 127449 77175 127759 85961
rect 127449 77147 127497 77175
rect 127525 77147 127559 77175
rect 127587 77147 127621 77175
rect 127649 77147 127683 77175
rect 127711 77147 127759 77175
rect 127449 77113 127759 77147
rect 127449 77085 127497 77113
rect 127525 77085 127559 77113
rect 127587 77085 127621 77113
rect 127649 77085 127683 77113
rect 127711 77085 127759 77113
rect 127449 77051 127759 77085
rect 127449 77023 127497 77051
rect 127525 77023 127559 77051
rect 127587 77023 127621 77051
rect 127649 77023 127683 77051
rect 127711 77023 127759 77051
rect 127449 76989 127759 77023
rect 127449 76961 127497 76989
rect 127525 76961 127559 76989
rect 127587 76961 127621 76989
rect 127649 76961 127683 76989
rect 127711 76961 127759 76989
rect 127449 68175 127759 76961
rect 127449 68147 127497 68175
rect 127525 68147 127559 68175
rect 127587 68147 127621 68175
rect 127649 68147 127683 68175
rect 127711 68147 127759 68175
rect 127449 68113 127759 68147
rect 127449 68085 127497 68113
rect 127525 68085 127559 68113
rect 127587 68085 127621 68113
rect 127649 68085 127683 68113
rect 127711 68085 127759 68113
rect 127449 68051 127759 68085
rect 127449 68023 127497 68051
rect 127525 68023 127559 68051
rect 127587 68023 127621 68051
rect 127649 68023 127683 68051
rect 127711 68023 127759 68051
rect 127449 67989 127759 68023
rect 127449 67961 127497 67989
rect 127525 67961 127559 67989
rect 127587 67961 127621 67989
rect 127649 67961 127683 67989
rect 127711 67961 127759 67989
rect 127449 59175 127759 67961
rect 127449 59147 127497 59175
rect 127525 59147 127559 59175
rect 127587 59147 127621 59175
rect 127649 59147 127683 59175
rect 127711 59147 127759 59175
rect 127449 59113 127759 59147
rect 127449 59085 127497 59113
rect 127525 59085 127559 59113
rect 127587 59085 127621 59113
rect 127649 59085 127683 59113
rect 127711 59085 127759 59113
rect 127449 59051 127759 59085
rect 127449 59023 127497 59051
rect 127525 59023 127559 59051
rect 127587 59023 127621 59051
rect 127649 59023 127683 59051
rect 127711 59023 127759 59051
rect 127449 58989 127759 59023
rect 127449 58961 127497 58989
rect 127525 58961 127559 58989
rect 127587 58961 127621 58989
rect 127649 58961 127683 58989
rect 127711 58961 127759 58989
rect 127449 50175 127759 58961
rect 127449 50147 127497 50175
rect 127525 50147 127559 50175
rect 127587 50147 127621 50175
rect 127649 50147 127683 50175
rect 127711 50147 127759 50175
rect 127449 50113 127759 50147
rect 127449 50085 127497 50113
rect 127525 50085 127559 50113
rect 127587 50085 127621 50113
rect 127649 50085 127683 50113
rect 127711 50085 127759 50113
rect 127449 50051 127759 50085
rect 127449 50023 127497 50051
rect 127525 50023 127559 50051
rect 127587 50023 127621 50051
rect 127649 50023 127683 50051
rect 127711 50023 127759 50051
rect 127449 49989 127759 50023
rect 127449 49961 127497 49989
rect 127525 49961 127559 49989
rect 127587 49961 127621 49989
rect 127649 49961 127683 49989
rect 127711 49961 127759 49989
rect 127449 41175 127759 49961
rect 127449 41147 127497 41175
rect 127525 41147 127559 41175
rect 127587 41147 127621 41175
rect 127649 41147 127683 41175
rect 127711 41147 127759 41175
rect 127449 41113 127759 41147
rect 127449 41085 127497 41113
rect 127525 41085 127559 41113
rect 127587 41085 127621 41113
rect 127649 41085 127683 41113
rect 127711 41085 127759 41113
rect 127449 41051 127759 41085
rect 127449 41023 127497 41051
rect 127525 41023 127559 41051
rect 127587 41023 127621 41051
rect 127649 41023 127683 41051
rect 127711 41023 127759 41051
rect 127449 40989 127759 41023
rect 127449 40961 127497 40989
rect 127525 40961 127559 40989
rect 127587 40961 127621 40989
rect 127649 40961 127683 40989
rect 127711 40961 127759 40989
rect 127449 32175 127759 40961
rect 127449 32147 127497 32175
rect 127525 32147 127559 32175
rect 127587 32147 127621 32175
rect 127649 32147 127683 32175
rect 127711 32147 127759 32175
rect 127449 32113 127759 32147
rect 127449 32085 127497 32113
rect 127525 32085 127559 32113
rect 127587 32085 127621 32113
rect 127649 32085 127683 32113
rect 127711 32085 127759 32113
rect 127449 32051 127759 32085
rect 127449 32023 127497 32051
rect 127525 32023 127559 32051
rect 127587 32023 127621 32051
rect 127649 32023 127683 32051
rect 127711 32023 127759 32051
rect 127449 31989 127759 32023
rect 127449 31961 127497 31989
rect 127525 31961 127559 31989
rect 127587 31961 127621 31989
rect 127649 31961 127683 31989
rect 127711 31961 127759 31989
rect 127449 23175 127759 31961
rect 127449 23147 127497 23175
rect 127525 23147 127559 23175
rect 127587 23147 127621 23175
rect 127649 23147 127683 23175
rect 127711 23147 127759 23175
rect 127449 23113 127759 23147
rect 127449 23085 127497 23113
rect 127525 23085 127559 23113
rect 127587 23085 127621 23113
rect 127649 23085 127683 23113
rect 127711 23085 127759 23113
rect 127449 23051 127759 23085
rect 127449 23023 127497 23051
rect 127525 23023 127559 23051
rect 127587 23023 127621 23051
rect 127649 23023 127683 23051
rect 127711 23023 127759 23051
rect 127449 22989 127759 23023
rect 127449 22961 127497 22989
rect 127525 22961 127559 22989
rect 127587 22961 127621 22989
rect 127649 22961 127683 22989
rect 127711 22961 127759 22989
rect 127449 14175 127759 22961
rect 127449 14147 127497 14175
rect 127525 14147 127559 14175
rect 127587 14147 127621 14175
rect 127649 14147 127683 14175
rect 127711 14147 127759 14175
rect 127449 14113 127759 14147
rect 127449 14085 127497 14113
rect 127525 14085 127559 14113
rect 127587 14085 127621 14113
rect 127649 14085 127683 14113
rect 127711 14085 127759 14113
rect 127449 14051 127759 14085
rect 127449 14023 127497 14051
rect 127525 14023 127559 14051
rect 127587 14023 127621 14051
rect 127649 14023 127683 14051
rect 127711 14023 127759 14051
rect 127449 13989 127759 14023
rect 127449 13961 127497 13989
rect 127525 13961 127559 13989
rect 127587 13961 127621 13989
rect 127649 13961 127683 13989
rect 127711 13961 127759 13989
rect 127449 5175 127759 13961
rect 127449 5147 127497 5175
rect 127525 5147 127559 5175
rect 127587 5147 127621 5175
rect 127649 5147 127683 5175
rect 127711 5147 127759 5175
rect 127449 5113 127759 5147
rect 127449 5085 127497 5113
rect 127525 5085 127559 5113
rect 127587 5085 127621 5113
rect 127649 5085 127683 5113
rect 127711 5085 127759 5113
rect 127449 5051 127759 5085
rect 127449 5023 127497 5051
rect 127525 5023 127559 5051
rect 127587 5023 127621 5051
rect 127649 5023 127683 5051
rect 127711 5023 127759 5051
rect 127449 4989 127759 5023
rect 127449 4961 127497 4989
rect 127525 4961 127559 4989
rect 127587 4961 127621 4989
rect 127649 4961 127683 4989
rect 127711 4961 127759 4989
rect 127449 -560 127759 4961
rect 127449 -588 127497 -560
rect 127525 -588 127559 -560
rect 127587 -588 127621 -560
rect 127649 -588 127683 -560
rect 127711 -588 127759 -560
rect 127449 -622 127759 -588
rect 127449 -650 127497 -622
rect 127525 -650 127559 -622
rect 127587 -650 127621 -622
rect 127649 -650 127683 -622
rect 127711 -650 127759 -622
rect 127449 -684 127759 -650
rect 127449 -712 127497 -684
rect 127525 -712 127559 -684
rect 127587 -712 127621 -684
rect 127649 -712 127683 -684
rect 127711 -712 127759 -684
rect 127449 -746 127759 -712
rect 127449 -774 127497 -746
rect 127525 -774 127559 -746
rect 127587 -774 127621 -746
rect 127649 -774 127683 -746
rect 127711 -774 127759 -746
rect 127449 -822 127759 -774
rect 140949 128175 141259 131025
rect 140949 128147 140997 128175
rect 141025 128147 141059 128175
rect 141087 128147 141121 128175
rect 141149 128147 141183 128175
rect 141211 128147 141259 128175
rect 140949 128113 141259 128147
rect 140949 128085 140997 128113
rect 141025 128085 141059 128113
rect 141087 128085 141121 128113
rect 141149 128085 141183 128113
rect 141211 128085 141259 128113
rect 140949 128051 141259 128085
rect 140949 128023 140997 128051
rect 141025 128023 141059 128051
rect 141087 128023 141121 128051
rect 141149 128023 141183 128051
rect 141211 128023 141259 128051
rect 140949 127989 141259 128023
rect 140949 127961 140997 127989
rect 141025 127961 141059 127989
rect 141087 127961 141121 127989
rect 141149 127961 141183 127989
rect 141211 127961 141259 127989
rect 140949 119175 141259 127961
rect 140949 119147 140997 119175
rect 141025 119147 141059 119175
rect 141087 119147 141121 119175
rect 141149 119147 141183 119175
rect 141211 119147 141259 119175
rect 140949 119113 141259 119147
rect 140949 119085 140997 119113
rect 141025 119085 141059 119113
rect 141087 119085 141121 119113
rect 141149 119085 141183 119113
rect 141211 119085 141259 119113
rect 140949 119051 141259 119085
rect 140949 119023 140997 119051
rect 141025 119023 141059 119051
rect 141087 119023 141121 119051
rect 141149 119023 141183 119051
rect 141211 119023 141259 119051
rect 140949 118989 141259 119023
rect 140949 118961 140997 118989
rect 141025 118961 141059 118989
rect 141087 118961 141121 118989
rect 141149 118961 141183 118989
rect 141211 118961 141259 118989
rect 140949 110175 141259 118961
rect 140949 110147 140997 110175
rect 141025 110147 141059 110175
rect 141087 110147 141121 110175
rect 141149 110147 141183 110175
rect 141211 110147 141259 110175
rect 140949 110113 141259 110147
rect 140949 110085 140997 110113
rect 141025 110085 141059 110113
rect 141087 110085 141121 110113
rect 141149 110085 141183 110113
rect 141211 110085 141259 110113
rect 140949 110051 141259 110085
rect 140949 110023 140997 110051
rect 141025 110023 141059 110051
rect 141087 110023 141121 110051
rect 141149 110023 141183 110051
rect 141211 110023 141259 110051
rect 140949 109989 141259 110023
rect 140949 109961 140997 109989
rect 141025 109961 141059 109989
rect 141087 109961 141121 109989
rect 141149 109961 141183 109989
rect 141211 109961 141259 109989
rect 140949 101175 141259 109961
rect 140949 101147 140997 101175
rect 141025 101147 141059 101175
rect 141087 101147 141121 101175
rect 141149 101147 141183 101175
rect 141211 101147 141259 101175
rect 140949 101113 141259 101147
rect 140949 101085 140997 101113
rect 141025 101085 141059 101113
rect 141087 101085 141121 101113
rect 141149 101085 141183 101113
rect 141211 101085 141259 101113
rect 140949 101051 141259 101085
rect 140949 101023 140997 101051
rect 141025 101023 141059 101051
rect 141087 101023 141121 101051
rect 141149 101023 141183 101051
rect 141211 101023 141259 101051
rect 140949 100989 141259 101023
rect 140949 100961 140997 100989
rect 141025 100961 141059 100989
rect 141087 100961 141121 100989
rect 141149 100961 141183 100989
rect 141211 100961 141259 100989
rect 140949 92175 141259 100961
rect 140949 92147 140997 92175
rect 141025 92147 141059 92175
rect 141087 92147 141121 92175
rect 141149 92147 141183 92175
rect 141211 92147 141259 92175
rect 140949 92113 141259 92147
rect 140949 92085 140997 92113
rect 141025 92085 141059 92113
rect 141087 92085 141121 92113
rect 141149 92085 141183 92113
rect 141211 92085 141259 92113
rect 140949 92051 141259 92085
rect 140949 92023 140997 92051
rect 141025 92023 141059 92051
rect 141087 92023 141121 92051
rect 141149 92023 141183 92051
rect 141211 92023 141259 92051
rect 140949 91989 141259 92023
rect 140949 91961 140997 91989
rect 141025 91961 141059 91989
rect 141087 91961 141121 91989
rect 141149 91961 141183 91989
rect 141211 91961 141259 91989
rect 140949 83175 141259 91961
rect 140949 83147 140997 83175
rect 141025 83147 141059 83175
rect 141087 83147 141121 83175
rect 141149 83147 141183 83175
rect 141211 83147 141259 83175
rect 140949 83113 141259 83147
rect 140949 83085 140997 83113
rect 141025 83085 141059 83113
rect 141087 83085 141121 83113
rect 141149 83085 141183 83113
rect 141211 83085 141259 83113
rect 140949 83051 141259 83085
rect 140949 83023 140997 83051
rect 141025 83023 141059 83051
rect 141087 83023 141121 83051
rect 141149 83023 141183 83051
rect 141211 83023 141259 83051
rect 140949 82989 141259 83023
rect 140949 82961 140997 82989
rect 141025 82961 141059 82989
rect 141087 82961 141121 82989
rect 141149 82961 141183 82989
rect 141211 82961 141259 82989
rect 140949 74175 141259 82961
rect 140949 74147 140997 74175
rect 141025 74147 141059 74175
rect 141087 74147 141121 74175
rect 141149 74147 141183 74175
rect 141211 74147 141259 74175
rect 140949 74113 141259 74147
rect 140949 74085 140997 74113
rect 141025 74085 141059 74113
rect 141087 74085 141121 74113
rect 141149 74085 141183 74113
rect 141211 74085 141259 74113
rect 140949 74051 141259 74085
rect 140949 74023 140997 74051
rect 141025 74023 141059 74051
rect 141087 74023 141121 74051
rect 141149 74023 141183 74051
rect 141211 74023 141259 74051
rect 140949 73989 141259 74023
rect 140949 73961 140997 73989
rect 141025 73961 141059 73989
rect 141087 73961 141121 73989
rect 141149 73961 141183 73989
rect 141211 73961 141259 73989
rect 140949 65175 141259 73961
rect 140949 65147 140997 65175
rect 141025 65147 141059 65175
rect 141087 65147 141121 65175
rect 141149 65147 141183 65175
rect 141211 65147 141259 65175
rect 140949 65113 141259 65147
rect 140949 65085 140997 65113
rect 141025 65085 141059 65113
rect 141087 65085 141121 65113
rect 141149 65085 141183 65113
rect 141211 65085 141259 65113
rect 140949 65051 141259 65085
rect 140949 65023 140997 65051
rect 141025 65023 141059 65051
rect 141087 65023 141121 65051
rect 141149 65023 141183 65051
rect 141211 65023 141259 65051
rect 140949 64989 141259 65023
rect 140949 64961 140997 64989
rect 141025 64961 141059 64989
rect 141087 64961 141121 64989
rect 141149 64961 141183 64989
rect 141211 64961 141259 64989
rect 140949 56175 141259 64961
rect 140949 56147 140997 56175
rect 141025 56147 141059 56175
rect 141087 56147 141121 56175
rect 141149 56147 141183 56175
rect 141211 56147 141259 56175
rect 140949 56113 141259 56147
rect 140949 56085 140997 56113
rect 141025 56085 141059 56113
rect 141087 56085 141121 56113
rect 141149 56085 141183 56113
rect 141211 56085 141259 56113
rect 140949 56051 141259 56085
rect 140949 56023 140997 56051
rect 141025 56023 141059 56051
rect 141087 56023 141121 56051
rect 141149 56023 141183 56051
rect 141211 56023 141259 56051
rect 140949 55989 141259 56023
rect 140949 55961 140997 55989
rect 141025 55961 141059 55989
rect 141087 55961 141121 55989
rect 141149 55961 141183 55989
rect 141211 55961 141259 55989
rect 140949 47175 141259 55961
rect 140949 47147 140997 47175
rect 141025 47147 141059 47175
rect 141087 47147 141121 47175
rect 141149 47147 141183 47175
rect 141211 47147 141259 47175
rect 140949 47113 141259 47147
rect 140949 47085 140997 47113
rect 141025 47085 141059 47113
rect 141087 47085 141121 47113
rect 141149 47085 141183 47113
rect 141211 47085 141259 47113
rect 140949 47051 141259 47085
rect 140949 47023 140997 47051
rect 141025 47023 141059 47051
rect 141087 47023 141121 47051
rect 141149 47023 141183 47051
rect 141211 47023 141259 47051
rect 140949 46989 141259 47023
rect 140949 46961 140997 46989
rect 141025 46961 141059 46989
rect 141087 46961 141121 46989
rect 141149 46961 141183 46989
rect 141211 46961 141259 46989
rect 140949 38175 141259 46961
rect 140949 38147 140997 38175
rect 141025 38147 141059 38175
rect 141087 38147 141121 38175
rect 141149 38147 141183 38175
rect 141211 38147 141259 38175
rect 140949 38113 141259 38147
rect 140949 38085 140997 38113
rect 141025 38085 141059 38113
rect 141087 38085 141121 38113
rect 141149 38085 141183 38113
rect 141211 38085 141259 38113
rect 140949 38051 141259 38085
rect 140949 38023 140997 38051
rect 141025 38023 141059 38051
rect 141087 38023 141121 38051
rect 141149 38023 141183 38051
rect 141211 38023 141259 38051
rect 140949 37989 141259 38023
rect 140949 37961 140997 37989
rect 141025 37961 141059 37989
rect 141087 37961 141121 37989
rect 141149 37961 141183 37989
rect 141211 37961 141259 37989
rect 140949 29175 141259 37961
rect 140949 29147 140997 29175
rect 141025 29147 141059 29175
rect 141087 29147 141121 29175
rect 141149 29147 141183 29175
rect 141211 29147 141259 29175
rect 140949 29113 141259 29147
rect 140949 29085 140997 29113
rect 141025 29085 141059 29113
rect 141087 29085 141121 29113
rect 141149 29085 141183 29113
rect 141211 29085 141259 29113
rect 140949 29051 141259 29085
rect 140949 29023 140997 29051
rect 141025 29023 141059 29051
rect 141087 29023 141121 29051
rect 141149 29023 141183 29051
rect 141211 29023 141259 29051
rect 140949 28989 141259 29023
rect 140949 28961 140997 28989
rect 141025 28961 141059 28989
rect 141087 28961 141121 28989
rect 141149 28961 141183 28989
rect 141211 28961 141259 28989
rect 140949 20175 141259 28961
rect 140949 20147 140997 20175
rect 141025 20147 141059 20175
rect 141087 20147 141121 20175
rect 141149 20147 141183 20175
rect 141211 20147 141259 20175
rect 140949 20113 141259 20147
rect 140949 20085 140997 20113
rect 141025 20085 141059 20113
rect 141087 20085 141121 20113
rect 141149 20085 141183 20113
rect 141211 20085 141259 20113
rect 140949 20051 141259 20085
rect 140949 20023 140997 20051
rect 141025 20023 141059 20051
rect 141087 20023 141121 20051
rect 141149 20023 141183 20051
rect 141211 20023 141259 20051
rect 140949 19989 141259 20023
rect 140949 19961 140997 19989
rect 141025 19961 141059 19989
rect 141087 19961 141121 19989
rect 141149 19961 141183 19989
rect 141211 19961 141259 19989
rect 140949 11175 141259 19961
rect 140949 11147 140997 11175
rect 141025 11147 141059 11175
rect 141087 11147 141121 11175
rect 141149 11147 141183 11175
rect 141211 11147 141259 11175
rect 140949 11113 141259 11147
rect 140949 11085 140997 11113
rect 141025 11085 141059 11113
rect 141087 11085 141121 11113
rect 141149 11085 141183 11113
rect 141211 11085 141259 11113
rect 140949 11051 141259 11085
rect 140949 11023 140997 11051
rect 141025 11023 141059 11051
rect 141087 11023 141121 11051
rect 141149 11023 141183 11051
rect 141211 11023 141259 11051
rect 140949 10989 141259 11023
rect 140949 10961 140997 10989
rect 141025 10961 141059 10989
rect 141087 10961 141121 10989
rect 141149 10961 141183 10989
rect 141211 10961 141259 10989
rect 140949 2175 141259 10961
rect 140949 2147 140997 2175
rect 141025 2147 141059 2175
rect 141087 2147 141121 2175
rect 141149 2147 141183 2175
rect 141211 2147 141259 2175
rect 140949 2113 141259 2147
rect 140949 2085 140997 2113
rect 141025 2085 141059 2113
rect 141087 2085 141121 2113
rect 141149 2085 141183 2113
rect 141211 2085 141259 2113
rect 140949 2051 141259 2085
rect 140949 2023 140997 2051
rect 141025 2023 141059 2051
rect 141087 2023 141121 2051
rect 141149 2023 141183 2051
rect 141211 2023 141259 2051
rect 140949 1989 141259 2023
rect 140949 1961 140997 1989
rect 141025 1961 141059 1989
rect 141087 1961 141121 1989
rect 141149 1961 141183 1989
rect 141211 1961 141259 1989
rect 140949 -80 141259 1961
rect 140949 -108 140997 -80
rect 141025 -108 141059 -80
rect 141087 -108 141121 -80
rect 141149 -108 141183 -80
rect 141211 -108 141259 -80
rect 140949 -142 141259 -108
rect 140949 -170 140997 -142
rect 141025 -170 141059 -142
rect 141087 -170 141121 -142
rect 141149 -170 141183 -142
rect 141211 -170 141259 -142
rect 140949 -204 141259 -170
rect 140949 -232 140997 -204
rect 141025 -232 141059 -204
rect 141087 -232 141121 -204
rect 141149 -232 141183 -204
rect 141211 -232 141259 -204
rect 140949 -266 141259 -232
rect 140949 -294 140997 -266
rect 141025 -294 141059 -266
rect 141087 -294 141121 -266
rect 141149 -294 141183 -266
rect 141211 -294 141259 -266
rect 140949 -822 141259 -294
rect 142809 131014 143119 131025
rect 142809 130986 142857 131014
rect 142885 130986 142919 131014
rect 142947 130986 142981 131014
rect 143009 130986 143043 131014
rect 143071 130986 143119 131014
rect 142809 130952 143119 130986
rect 142809 130924 142857 130952
rect 142885 130924 142919 130952
rect 142947 130924 142981 130952
rect 143009 130924 143043 130952
rect 143071 130924 143119 130952
rect 142809 122175 143119 130924
rect 142809 122147 142857 122175
rect 142885 122147 142919 122175
rect 142947 122147 142981 122175
rect 143009 122147 143043 122175
rect 143071 122147 143119 122175
rect 142809 122113 143119 122147
rect 142809 122085 142857 122113
rect 142885 122085 142919 122113
rect 142947 122085 142981 122113
rect 143009 122085 143043 122113
rect 143071 122085 143119 122113
rect 142809 122051 143119 122085
rect 142809 122023 142857 122051
rect 142885 122023 142919 122051
rect 142947 122023 142981 122051
rect 143009 122023 143043 122051
rect 143071 122023 143119 122051
rect 142809 121989 143119 122023
rect 142809 121961 142857 121989
rect 142885 121961 142919 121989
rect 142947 121961 142981 121989
rect 143009 121961 143043 121989
rect 143071 121961 143119 121989
rect 142809 113175 143119 121961
rect 142809 113147 142857 113175
rect 142885 113147 142919 113175
rect 142947 113147 142981 113175
rect 143009 113147 143043 113175
rect 143071 113147 143119 113175
rect 142809 113113 143119 113147
rect 142809 113085 142857 113113
rect 142885 113085 142919 113113
rect 142947 113085 142981 113113
rect 143009 113085 143043 113113
rect 143071 113085 143119 113113
rect 142809 113051 143119 113085
rect 142809 113023 142857 113051
rect 142885 113023 142919 113051
rect 142947 113023 142981 113051
rect 143009 113023 143043 113051
rect 143071 113023 143119 113051
rect 142809 112989 143119 113023
rect 142809 112961 142857 112989
rect 142885 112961 142919 112989
rect 142947 112961 142981 112989
rect 143009 112961 143043 112989
rect 143071 112961 143119 112989
rect 142809 104175 143119 112961
rect 142809 104147 142857 104175
rect 142885 104147 142919 104175
rect 142947 104147 142981 104175
rect 143009 104147 143043 104175
rect 143071 104147 143119 104175
rect 142809 104113 143119 104147
rect 142809 104085 142857 104113
rect 142885 104085 142919 104113
rect 142947 104085 142981 104113
rect 143009 104085 143043 104113
rect 143071 104085 143119 104113
rect 142809 104051 143119 104085
rect 142809 104023 142857 104051
rect 142885 104023 142919 104051
rect 142947 104023 142981 104051
rect 143009 104023 143043 104051
rect 143071 104023 143119 104051
rect 142809 103989 143119 104023
rect 142809 103961 142857 103989
rect 142885 103961 142919 103989
rect 142947 103961 142981 103989
rect 143009 103961 143043 103989
rect 143071 103961 143119 103989
rect 142809 95175 143119 103961
rect 142809 95147 142857 95175
rect 142885 95147 142919 95175
rect 142947 95147 142981 95175
rect 143009 95147 143043 95175
rect 143071 95147 143119 95175
rect 142809 95113 143119 95147
rect 142809 95085 142857 95113
rect 142885 95085 142919 95113
rect 142947 95085 142981 95113
rect 143009 95085 143043 95113
rect 143071 95085 143119 95113
rect 142809 95051 143119 95085
rect 142809 95023 142857 95051
rect 142885 95023 142919 95051
rect 142947 95023 142981 95051
rect 143009 95023 143043 95051
rect 143071 95023 143119 95051
rect 142809 94989 143119 95023
rect 142809 94961 142857 94989
rect 142885 94961 142919 94989
rect 142947 94961 142981 94989
rect 143009 94961 143043 94989
rect 143071 94961 143119 94989
rect 142809 86175 143119 94961
rect 142809 86147 142857 86175
rect 142885 86147 142919 86175
rect 142947 86147 142981 86175
rect 143009 86147 143043 86175
rect 143071 86147 143119 86175
rect 142809 86113 143119 86147
rect 142809 86085 142857 86113
rect 142885 86085 142919 86113
rect 142947 86085 142981 86113
rect 143009 86085 143043 86113
rect 143071 86085 143119 86113
rect 142809 86051 143119 86085
rect 142809 86023 142857 86051
rect 142885 86023 142919 86051
rect 142947 86023 142981 86051
rect 143009 86023 143043 86051
rect 143071 86023 143119 86051
rect 142809 85989 143119 86023
rect 142809 85961 142857 85989
rect 142885 85961 142919 85989
rect 142947 85961 142981 85989
rect 143009 85961 143043 85989
rect 143071 85961 143119 85989
rect 142809 77175 143119 85961
rect 142809 77147 142857 77175
rect 142885 77147 142919 77175
rect 142947 77147 142981 77175
rect 143009 77147 143043 77175
rect 143071 77147 143119 77175
rect 142809 77113 143119 77147
rect 142809 77085 142857 77113
rect 142885 77085 142919 77113
rect 142947 77085 142981 77113
rect 143009 77085 143043 77113
rect 143071 77085 143119 77113
rect 142809 77051 143119 77085
rect 142809 77023 142857 77051
rect 142885 77023 142919 77051
rect 142947 77023 142981 77051
rect 143009 77023 143043 77051
rect 143071 77023 143119 77051
rect 142809 76989 143119 77023
rect 142809 76961 142857 76989
rect 142885 76961 142919 76989
rect 142947 76961 142981 76989
rect 143009 76961 143043 76989
rect 143071 76961 143119 76989
rect 142809 68175 143119 76961
rect 142809 68147 142857 68175
rect 142885 68147 142919 68175
rect 142947 68147 142981 68175
rect 143009 68147 143043 68175
rect 143071 68147 143119 68175
rect 142809 68113 143119 68147
rect 142809 68085 142857 68113
rect 142885 68085 142919 68113
rect 142947 68085 142981 68113
rect 143009 68085 143043 68113
rect 143071 68085 143119 68113
rect 142809 68051 143119 68085
rect 142809 68023 142857 68051
rect 142885 68023 142919 68051
rect 142947 68023 142981 68051
rect 143009 68023 143043 68051
rect 143071 68023 143119 68051
rect 142809 67989 143119 68023
rect 142809 67961 142857 67989
rect 142885 67961 142919 67989
rect 142947 67961 142981 67989
rect 143009 67961 143043 67989
rect 143071 67961 143119 67989
rect 142809 59175 143119 67961
rect 142809 59147 142857 59175
rect 142885 59147 142919 59175
rect 142947 59147 142981 59175
rect 143009 59147 143043 59175
rect 143071 59147 143119 59175
rect 142809 59113 143119 59147
rect 142809 59085 142857 59113
rect 142885 59085 142919 59113
rect 142947 59085 142981 59113
rect 143009 59085 143043 59113
rect 143071 59085 143119 59113
rect 142809 59051 143119 59085
rect 142809 59023 142857 59051
rect 142885 59023 142919 59051
rect 142947 59023 142981 59051
rect 143009 59023 143043 59051
rect 143071 59023 143119 59051
rect 142809 58989 143119 59023
rect 142809 58961 142857 58989
rect 142885 58961 142919 58989
rect 142947 58961 142981 58989
rect 143009 58961 143043 58989
rect 143071 58961 143119 58989
rect 142809 50175 143119 58961
rect 142809 50147 142857 50175
rect 142885 50147 142919 50175
rect 142947 50147 142981 50175
rect 143009 50147 143043 50175
rect 143071 50147 143119 50175
rect 142809 50113 143119 50147
rect 142809 50085 142857 50113
rect 142885 50085 142919 50113
rect 142947 50085 142981 50113
rect 143009 50085 143043 50113
rect 143071 50085 143119 50113
rect 142809 50051 143119 50085
rect 142809 50023 142857 50051
rect 142885 50023 142919 50051
rect 142947 50023 142981 50051
rect 143009 50023 143043 50051
rect 143071 50023 143119 50051
rect 142809 49989 143119 50023
rect 142809 49961 142857 49989
rect 142885 49961 142919 49989
rect 142947 49961 142981 49989
rect 143009 49961 143043 49989
rect 143071 49961 143119 49989
rect 142809 41175 143119 49961
rect 142809 41147 142857 41175
rect 142885 41147 142919 41175
rect 142947 41147 142981 41175
rect 143009 41147 143043 41175
rect 143071 41147 143119 41175
rect 142809 41113 143119 41147
rect 142809 41085 142857 41113
rect 142885 41085 142919 41113
rect 142947 41085 142981 41113
rect 143009 41085 143043 41113
rect 143071 41085 143119 41113
rect 142809 41051 143119 41085
rect 142809 41023 142857 41051
rect 142885 41023 142919 41051
rect 142947 41023 142981 41051
rect 143009 41023 143043 41051
rect 143071 41023 143119 41051
rect 142809 40989 143119 41023
rect 142809 40961 142857 40989
rect 142885 40961 142919 40989
rect 142947 40961 142981 40989
rect 143009 40961 143043 40989
rect 143071 40961 143119 40989
rect 142809 32175 143119 40961
rect 142809 32147 142857 32175
rect 142885 32147 142919 32175
rect 142947 32147 142981 32175
rect 143009 32147 143043 32175
rect 143071 32147 143119 32175
rect 142809 32113 143119 32147
rect 142809 32085 142857 32113
rect 142885 32085 142919 32113
rect 142947 32085 142981 32113
rect 143009 32085 143043 32113
rect 143071 32085 143119 32113
rect 142809 32051 143119 32085
rect 142809 32023 142857 32051
rect 142885 32023 142919 32051
rect 142947 32023 142981 32051
rect 143009 32023 143043 32051
rect 143071 32023 143119 32051
rect 142809 31989 143119 32023
rect 142809 31961 142857 31989
rect 142885 31961 142919 31989
rect 142947 31961 142981 31989
rect 143009 31961 143043 31989
rect 143071 31961 143119 31989
rect 142809 23175 143119 31961
rect 142809 23147 142857 23175
rect 142885 23147 142919 23175
rect 142947 23147 142981 23175
rect 143009 23147 143043 23175
rect 143071 23147 143119 23175
rect 142809 23113 143119 23147
rect 142809 23085 142857 23113
rect 142885 23085 142919 23113
rect 142947 23085 142981 23113
rect 143009 23085 143043 23113
rect 143071 23085 143119 23113
rect 142809 23051 143119 23085
rect 142809 23023 142857 23051
rect 142885 23023 142919 23051
rect 142947 23023 142981 23051
rect 143009 23023 143043 23051
rect 143071 23023 143119 23051
rect 142809 22989 143119 23023
rect 142809 22961 142857 22989
rect 142885 22961 142919 22989
rect 142947 22961 142981 22989
rect 143009 22961 143043 22989
rect 143071 22961 143119 22989
rect 142809 14175 143119 22961
rect 142809 14147 142857 14175
rect 142885 14147 142919 14175
rect 142947 14147 142981 14175
rect 143009 14147 143043 14175
rect 143071 14147 143119 14175
rect 142809 14113 143119 14147
rect 142809 14085 142857 14113
rect 142885 14085 142919 14113
rect 142947 14085 142981 14113
rect 143009 14085 143043 14113
rect 143071 14085 143119 14113
rect 142809 14051 143119 14085
rect 142809 14023 142857 14051
rect 142885 14023 142919 14051
rect 142947 14023 142981 14051
rect 143009 14023 143043 14051
rect 143071 14023 143119 14051
rect 142809 13989 143119 14023
rect 142809 13961 142857 13989
rect 142885 13961 142919 13989
rect 142947 13961 142981 13989
rect 143009 13961 143043 13989
rect 143071 13961 143119 13989
rect 142809 5175 143119 13961
rect 142809 5147 142857 5175
rect 142885 5147 142919 5175
rect 142947 5147 142981 5175
rect 143009 5147 143043 5175
rect 143071 5147 143119 5175
rect 142809 5113 143119 5147
rect 142809 5085 142857 5113
rect 142885 5085 142919 5113
rect 142947 5085 142981 5113
rect 143009 5085 143043 5113
rect 143071 5085 143119 5113
rect 142809 5051 143119 5085
rect 142809 5023 142857 5051
rect 142885 5023 142919 5051
rect 142947 5023 142981 5051
rect 143009 5023 143043 5051
rect 143071 5023 143119 5051
rect 142809 4989 143119 5023
rect 142809 4961 142857 4989
rect 142885 4961 142919 4989
rect 142947 4961 142981 4989
rect 143009 4961 143043 4989
rect 143071 4961 143119 4989
rect 142809 -560 143119 4961
rect 142809 -588 142857 -560
rect 142885 -588 142919 -560
rect 142947 -588 142981 -560
rect 143009 -588 143043 -560
rect 143071 -588 143119 -560
rect 142809 -622 143119 -588
rect 142809 -650 142857 -622
rect 142885 -650 142919 -622
rect 142947 -650 142981 -622
rect 143009 -650 143043 -622
rect 143071 -650 143119 -622
rect 142809 -684 143119 -650
rect 142809 -712 142857 -684
rect 142885 -712 142919 -684
rect 142947 -712 142981 -684
rect 143009 -712 143043 -684
rect 143071 -712 143119 -684
rect 142809 -746 143119 -712
rect 142809 -774 142857 -746
rect 142885 -774 142919 -746
rect 142947 -774 142981 -746
rect 143009 -774 143043 -746
rect 143071 -774 143119 -746
rect 142809 -822 143119 -774
rect 156309 128175 156619 131025
rect 156309 128147 156357 128175
rect 156385 128147 156419 128175
rect 156447 128147 156481 128175
rect 156509 128147 156543 128175
rect 156571 128147 156619 128175
rect 156309 128113 156619 128147
rect 156309 128085 156357 128113
rect 156385 128085 156419 128113
rect 156447 128085 156481 128113
rect 156509 128085 156543 128113
rect 156571 128085 156619 128113
rect 156309 128051 156619 128085
rect 156309 128023 156357 128051
rect 156385 128023 156419 128051
rect 156447 128023 156481 128051
rect 156509 128023 156543 128051
rect 156571 128023 156619 128051
rect 156309 127989 156619 128023
rect 156309 127961 156357 127989
rect 156385 127961 156419 127989
rect 156447 127961 156481 127989
rect 156509 127961 156543 127989
rect 156571 127961 156619 127989
rect 156309 119175 156619 127961
rect 156309 119147 156357 119175
rect 156385 119147 156419 119175
rect 156447 119147 156481 119175
rect 156509 119147 156543 119175
rect 156571 119147 156619 119175
rect 156309 119113 156619 119147
rect 156309 119085 156357 119113
rect 156385 119085 156419 119113
rect 156447 119085 156481 119113
rect 156509 119085 156543 119113
rect 156571 119085 156619 119113
rect 156309 119051 156619 119085
rect 156309 119023 156357 119051
rect 156385 119023 156419 119051
rect 156447 119023 156481 119051
rect 156509 119023 156543 119051
rect 156571 119023 156619 119051
rect 156309 118989 156619 119023
rect 156309 118961 156357 118989
rect 156385 118961 156419 118989
rect 156447 118961 156481 118989
rect 156509 118961 156543 118989
rect 156571 118961 156619 118989
rect 156309 110175 156619 118961
rect 156309 110147 156357 110175
rect 156385 110147 156419 110175
rect 156447 110147 156481 110175
rect 156509 110147 156543 110175
rect 156571 110147 156619 110175
rect 156309 110113 156619 110147
rect 156309 110085 156357 110113
rect 156385 110085 156419 110113
rect 156447 110085 156481 110113
rect 156509 110085 156543 110113
rect 156571 110085 156619 110113
rect 156309 110051 156619 110085
rect 156309 110023 156357 110051
rect 156385 110023 156419 110051
rect 156447 110023 156481 110051
rect 156509 110023 156543 110051
rect 156571 110023 156619 110051
rect 156309 109989 156619 110023
rect 156309 109961 156357 109989
rect 156385 109961 156419 109989
rect 156447 109961 156481 109989
rect 156509 109961 156543 109989
rect 156571 109961 156619 109989
rect 156309 101175 156619 109961
rect 156309 101147 156357 101175
rect 156385 101147 156419 101175
rect 156447 101147 156481 101175
rect 156509 101147 156543 101175
rect 156571 101147 156619 101175
rect 156309 101113 156619 101147
rect 156309 101085 156357 101113
rect 156385 101085 156419 101113
rect 156447 101085 156481 101113
rect 156509 101085 156543 101113
rect 156571 101085 156619 101113
rect 156309 101051 156619 101085
rect 156309 101023 156357 101051
rect 156385 101023 156419 101051
rect 156447 101023 156481 101051
rect 156509 101023 156543 101051
rect 156571 101023 156619 101051
rect 156309 100989 156619 101023
rect 156309 100961 156357 100989
rect 156385 100961 156419 100989
rect 156447 100961 156481 100989
rect 156509 100961 156543 100989
rect 156571 100961 156619 100989
rect 156309 92175 156619 100961
rect 156309 92147 156357 92175
rect 156385 92147 156419 92175
rect 156447 92147 156481 92175
rect 156509 92147 156543 92175
rect 156571 92147 156619 92175
rect 156309 92113 156619 92147
rect 156309 92085 156357 92113
rect 156385 92085 156419 92113
rect 156447 92085 156481 92113
rect 156509 92085 156543 92113
rect 156571 92085 156619 92113
rect 156309 92051 156619 92085
rect 156309 92023 156357 92051
rect 156385 92023 156419 92051
rect 156447 92023 156481 92051
rect 156509 92023 156543 92051
rect 156571 92023 156619 92051
rect 156309 91989 156619 92023
rect 156309 91961 156357 91989
rect 156385 91961 156419 91989
rect 156447 91961 156481 91989
rect 156509 91961 156543 91989
rect 156571 91961 156619 91989
rect 156309 83175 156619 91961
rect 156309 83147 156357 83175
rect 156385 83147 156419 83175
rect 156447 83147 156481 83175
rect 156509 83147 156543 83175
rect 156571 83147 156619 83175
rect 156309 83113 156619 83147
rect 156309 83085 156357 83113
rect 156385 83085 156419 83113
rect 156447 83085 156481 83113
rect 156509 83085 156543 83113
rect 156571 83085 156619 83113
rect 156309 83051 156619 83085
rect 156309 83023 156357 83051
rect 156385 83023 156419 83051
rect 156447 83023 156481 83051
rect 156509 83023 156543 83051
rect 156571 83023 156619 83051
rect 156309 82989 156619 83023
rect 156309 82961 156357 82989
rect 156385 82961 156419 82989
rect 156447 82961 156481 82989
rect 156509 82961 156543 82989
rect 156571 82961 156619 82989
rect 156309 74175 156619 82961
rect 156309 74147 156357 74175
rect 156385 74147 156419 74175
rect 156447 74147 156481 74175
rect 156509 74147 156543 74175
rect 156571 74147 156619 74175
rect 156309 74113 156619 74147
rect 156309 74085 156357 74113
rect 156385 74085 156419 74113
rect 156447 74085 156481 74113
rect 156509 74085 156543 74113
rect 156571 74085 156619 74113
rect 156309 74051 156619 74085
rect 156309 74023 156357 74051
rect 156385 74023 156419 74051
rect 156447 74023 156481 74051
rect 156509 74023 156543 74051
rect 156571 74023 156619 74051
rect 156309 73989 156619 74023
rect 156309 73961 156357 73989
rect 156385 73961 156419 73989
rect 156447 73961 156481 73989
rect 156509 73961 156543 73989
rect 156571 73961 156619 73989
rect 156309 65175 156619 73961
rect 156309 65147 156357 65175
rect 156385 65147 156419 65175
rect 156447 65147 156481 65175
rect 156509 65147 156543 65175
rect 156571 65147 156619 65175
rect 156309 65113 156619 65147
rect 156309 65085 156357 65113
rect 156385 65085 156419 65113
rect 156447 65085 156481 65113
rect 156509 65085 156543 65113
rect 156571 65085 156619 65113
rect 156309 65051 156619 65085
rect 156309 65023 156357 65051
rect 156385 65023 156419 65051
rect 156447 65023 156481 65051
rect 156509 65023 156543 65051
rect 156571 65023 156619 65051
rect 156309 64989 156619 65023
rect 156309 64961 156357 64989
rect 156385 64961 156419 64989
rect 156447 64961 156481 64989
rect 156509 64961 156543 64989
rect 156571 64961 156619 64989
rect 156309 56175 156619 64961
rect 156309 56147 156357 56175
rect 156385 56147 156419 56175
rect 156447 56147 156481 56175
rect 156509 56147 156543 56175
rect 156571 56147 156619 56175
rect 156309 56113 156619 56147
rect 156309 56085 156357 56113
rect 156385 56085 156419 56113
rect 156447 56085 156481 56113
rect 156509 56085 156543 56113
rect 156571 56085 156619 56113
rect 156309 56051 156619 56085
rect 156309 56023 156357 56051
rect 156385 56023 156419 56051
rect 156447 56023 156481 56051
rect 156509 56023 156543 56051
rect 156571 56023 156619 56051
rect 156309 55989 156619 56023
rect 156309 55961 156357 55989
rect 156385 55961 156419 55989
rect 156447 55961 156481 55989
rect 156509 55961 156543 55989
rect 156571 55961 156619 55989
rect 156309 47175 156619 55961
rect 156309 47147 156357 47175
rect 156385 47147 156419 47175
rect 156447 47147 156481 47175
rect 156509 47147 156543 47175
rect 156571 47147 156619 47175
rect 156309 47113 156619 47147
rect 156309 47085 156357 47113
rect 156385 47085 156419 47113
rect 156447 47085 156481 47113
rect 156509 47085 156543 47113
rect 156571 47085 156619 47113
rect 156309 47051 156619 47085
rect 156309 47023 156357 47051
rect 156385 47023 156419 47051
rect 156447 47023 156481 47051
rect 156509 47023 156543 47051
rect 156571 47023 156619 47051
rect 156309 46989 156619 47023
rect 156309 46961 156357 46989
rect 156385 46961 156419 46989
rect 156447 46961 156481 46989
rect 156509 46961 156543 46989
rect 156571 46961 156619 46989
rect 156309 38175 156619 46961
rect 156309 38147 156357 38175
rect 156385 38147 156419 38175
rect 156447 38147 156481 38175
rect 156509 38147 156543 38175
rect 156571 38147 156619 38175
rect 156309 38113 156619 38147
rect 156309 38085 156357 38113
rect 156385 38085 156419 38113
rect 156447 38085 156481 38113
rect 156509 38085 156543 38113
rect 156571 38085 156619 38113
rect 156309 38051 156619 38085
rect 156309 38023 156357 38051
rect 156385 38023 156419 38051
rect 156447 38023 156481 38051
rect 156509 38023 156543 38051
rect 156571 38023 156619 38051
rect 156309 37989 156619 38023
rect 156309 37961 156357 37989
rect 156385 37961 156419 37989
rect 156447 37961 156481 37989
rect 156509 37961 156543 37989
rect 156571 37961 156619 37989
rect 156309 29175 156619 37961
rect 156309 29147 156357 29175
rect 156385 29147 156419 29175
rect 156447 29147 156481 29175
rect 156509 29147 156543 29175
rect 156571 29147 156619 29175
rect 156309 29113 156619 29147
rect 156309 29085 156357 29113
rect 156385 29085 156419 29113
rect 156447 29085 156481 29113
rect 156509 29085 156543 29113
rect 156571 29085 156619 29113
rect 156309 29051 156619 29085
rect 156309 29023 156357 29051
rect 156385 29023 156419 29051
rect 156447 29023 156481 29051
rect 156509 29023 156543 29051
rect 156571 29023 156619 29051
rect 156309 28989 156619 29023
rect 156309 28961 156357 28989
rect 156385 28961 156419 28989
rect 156447 28961 156481 28989
rect 156509 28961 156543 28989
rect 156571 28961 156619 28989
rect 156309 20175 156619 28961
rect 156309 20147 156357 20175
rect 156385 20147 156419 20175
rect 156447 20147 156481 20175
rect 156509 20147 156543 20175
rect 156571 20147 156619 20175
rect 156309 20113 156619 20147
rect 156309 20085 156357 20113
rect 156385 20085 156419 20113
rect 156447 20085 156481 20113
rect 156509 20085 156543 20113
rect 156571 20085 156619 20113
rect 156309 20051 156619 20085
rect 156309 20023 156357 20051
rect 156385 20023 156419 20051
rect 156447 20023 156481 20051
rect 156509 20023 156543 20051
rect 156571 20023 156619 20051
rect 156309 19989 156619 20023
rect 156309 19961 156357 19989
rect 156385 19961 156419 19989
rect 156447 19961 156481 19989
rect 156509 19961 156543 19989
rect 156571 19961 156619 19989
rect 156309 11175 156619 19961
rect 156309 11147 156357 11175
rect 156385 11147 156419 11175
rect 156447 11147 156481 11175
rect 156509 11147 156543 11175
rect 156571 11147 156619 11175
rect 156309 11113 156619 11147
rect 156309 11085 156357 11113
rect 156385 11085 156419 11113
rect 156447 11085 156481 11113
rect 156509 11085 156543 11113
rect 156571 11085 156619 11113
rect 156309 11051 156619 11085
rect 156309 11023 156357 11051
rect 156385 11023 156419 11051
rect 156447 11023 156481 11051
rect 156509 11023 156543 11051
rect 156571 11023 156619 11051
rect 156309 10989 156619 11023
rect 156309 10961 156357 10989
rect 156385 10961 156419 10989
rect 156447 10961 156481 10989
rect 156509 10961 156543 10989
rect 156571 10961 156619 10989
rect 156309 2175 156619 10961
rect 156309 2147 156357 2175
rect 156385 2147 156419 2175
rect 156447 2147 156481 2175
rect 156509 2147 156543 2175
rect 156571 2147 156619 2175
rect 156309 2113 156619 2147
rect 156309 2085 156357 2113
rect 156385 2085 156419 2113
rect 156447 2085 156481 2113
rect 156509 2085 156543 2113
rect 156571 2085 156619 2113
rect 156309 2051 156619 2085
rect 156309 2023 156357 2051
rect 156385 2023 156419 2051
rect 156447 2023 156481 2051
rect 156509 2023 156543 2051
rect 156571 2023 156619 2051
rect 156309 1989 156619 2023
rect 156309 1961 156357 1989
rect 156385 1961 156419 1989
rect 156447 1961 156481 1989
rect 156509 1961 156543 1989
rect 156571 1961 156619 1989
rect 156309 -80 156619 1961
rect 156309 -108 156357 -80
rect 156385 -108 156419 -80
rect 156447 -108 156481 -80
rect 156509 -108 156543 -80
rect 156571 -108 156619 -80
rect 156309 -142 156619 -108
rect 156309 -170 156357 -142
rect 156385 -170 156419 -142
rect 156447 -170 156481 -142
rect 156509 -170 156543 -142
rect 156571 -170 156619 -142
rect 156309 -204 156619 -170
rect 156309 -232 156357 -204
rect 156385 -232 156419 -204
rect 156447 -232 156481 -204
rect 156509 -232 156543 -204
rect 156571 -232 156619 -204
rect 156309 -266 156619 -232
rect 156309 -294 156357 -266
rect 156385 -294 156419 -266
rect 156447 -294 156481 -266
rect 156509 -294 156543 -266
rect 156571 -294 156619 -266
rect 156309 -822 156619 -294
rect 158169 131014 158479 131025
rect 158169 130986 158217 131014
rect 158245 130986 158279 131014
rect 158307 130986 158341 131014
rect 158369 130986 158403 131014
rect 158431 130986 158479 131014
rect 158169 130952 158479 130986
rect 158169 130924 158217 130952
rect 158245 130924 158279 130952
rect 158307 130924 158341 130952
rect 158369 130924 158403 130952
rect 158431 130924 158479 130952
rect 158169 122175 158479 130924
rect 173529 131014 173839 131025
rect 173529 130986 173577 131014
rect 173605 130986 173639 131014
rect 173667 130986 173701 131014
rect 173729 130986 173763 131014
rect 173791 130986 173839 131014
rect 173529 130952 173839 130986
rect 173529 130924 173577 130952
rect 173605 130924 173639 130952
rect 173667 130924 173701 130952
rect 173729 130924 173763 130952
rect 173791 130924 173839 130952
rect 173529 125367 173839 130924
rect 188889 131014 189199 131025
rect 188889 130986 188937 131014
rect 188965 130986 188999 131014
rect 189027 130986 189061 131014
rect 189089 130986 189123 131014
rect 189151 130986 189199 131014
rect 188889 130952 189199 130986
rect 188889 130924 188937 130952
rect 188965 130924 188999 130952
rect 189027 130924 189061 130952
rect 189089 130924 189123 130952
rect 189151 130924 189199 130952
rect 188889 125367 189199 130924
rect 204249 131023 204297 131051
rect 204325 131023 204359 131051
rect 204387 131023 204421 131051
rect 204449 131023 204483 131051
rect 204511 131023 204559 131051
rect 204249 130989 204559 131023
rect 204249 130961 204297 130989
rect 204325 130961 204359 130989
rect 204387 130961 204421 130989
rect 204449 130961 204483 130989
rect 204511 130961 204559 130989
rect 204249 125367 204559 130961
rect 217749 128175 218059 136961
rect 217749 128147 217797 128175
rect 217825 128147 217859 128175
rect 217887 128147 217921 128175
rect 217949 128147 217983 128175
rect 218011 128147 218059 128175
rect 217749 128113 218059 128147
rect 217749 128085 217797 128113
rect 217825 128085 217859 128113
rect 217887 128085 217921 128113
rect 217949 128085 217983 128113
rect 218011 128085 218059 128113
rect 217749 128051 218059 128085
rect 217749 128023 217797 128051
rect 217825 128023 217859 128051
rect 217887 128023 217921 128051
rect 217949 128023 217983 128051
rect 218011 128023 218059 128051
rect 217749 127989 218059 128023
rect 217749 127961 217797 127989
rect 217825 127961 217859 127989
rect 217887 127961 217921 127989
rect 217949 127961 217983 127989
rect 218011 127961 218059 127989
rect 217749 125367 218059 127961
rect 219609 299086 219919 299134
rect 219609 299058 219657 299086
rect 219685 299058 219719 299086
rect 219747 299058 219781 299086
rect 219809 299058 219843 299086
rect 219871 299058 219919 299086
rect 219609 299024 219919 299058
rect 219609 298996 219657 299024
rect 219685 298996 219719 299024
rect 219747 298996 219781 299024
rect 219809 298996 219843 299024
rect 219871 298996 219919 299024
rect 219609 298962 219919 298996
rect 219609 298934 219657 298962
rect 219685 298934 219719 298962
rect 219747 298934 219781 298962
rect 219809 298934 219843 298962
rect 219871 298934 219919 298962
rect 219609 298900 219919 298934
rect 219609 298872 219657 298900
rect 219685 298872 219719 298900
rect 219747 298872 219781 298900
rect 219809 298872 219843 298900
rect 219871 298872 219919 298900
rect 219609 293175 219919 298872
rect 219609 293147 219657 293175
rect 219685 293147 219719 293175
rect 219747 293147 219781 293175
rect 219809 293147 219843 293175
rect 219871 293147 219919 293175
rect 219609 293113 219919 293147
rect 219609 293085 219657 293113
rect 219685 293085 219719 293113
rect 219747 293085 219781 293113
rect 219809 293085 219843 293113
rect 219871 293085 219919 293113
rect 219609 293051 219919 293085
rect 219609 293023 219657 293051
rect 219685 293023 219719 293051
rect 219747 293023 219781 293051
rect 219809 293023 219843 293051
rect 219871 293023 219919 293051
rect 219609 292989 219919 293023
rect 219609 292961 219657 292989
rect 219685 292961 219719 292989
rect 219747 292961 219781 292989
rect 219809 292961 219843 292989
rect 219871 292961 219919 292989
rect 219609 284175 219919 292961
rect 219609 284147 219657 284175
rect 219685 284147 219719 284175
rect 219747 284147 219781 284175
rect 219809 284147 219843 284175
rect 219871 284147 219919 284175
rect 219609 284113 219919 284147
rect 219609 284085 219657 284113
rect 219685 284085 219719 284113
rect 219747 284085 219781 284113
rect 219809 284085 219843 284113
rect 219871 284085 219919 284113
rect 219609 284051 219919 284085
rect 219609 284023 219657 284051
rect 219685 284023 219719 284051
rect 219747 284023 219781 284051
rect 219809 284023 219843 284051
rect 219871 284023 219919 284051
rect 219609 283989 219919 284023
rect 219609 283961 219657 283989
rect 219685 283961 219719 283989
rect 219747 283961 219781 283989
rect 219809 283961 219843 283989
rect 219871 283961 219919 283989
rect 219609 275175 219919 283961
rect 219609 275147 219657 275175
rect 219685 275147 219719 275175
rect 219747 275147 219781 275175
rect 219809 275147 219843 275175
rect 219871 275147 219919 275175
rect 219609 275113 219919 275147
rect 219609 275085 219657 275113
rect 219685 275085 219719 275113
rect 219747 275085 219781 275113
rect 219809 275085 219843 275113
rect 219871 275085 219919 275113
rect 219609 275051 219919 275085
rect 219609 275023 219657 275051
rect 219685 275023 219719 275051
rect 219747 275023 219781 275051
rect 219809 275023 219843 275051
rect 219871 275023 219919 275051
rect 219609 274989 219919 275023
rect 219609 274961 219657 274989
rect 219685 274961 219719 274989
rect 219747 274961 219781 274989
rect 219809 274961 219843 274989
rect 219871 274961 219919 274989
rect 219609 266175 219919 274961
rect 219609 266147 219657 266175
rect 219685 266147 219719 266175
rect 219747 266147 219781 266175
rect 219809 266147 219843 266175
rect 219871 266147 219919 266175
rect 219609 266113 219919 266147
rect 219609 266085 219657 266113
rect 219685 266085 219719 266113
rect 219747 266085 219781 266113
rect 219809 266085 219843 266113
rect 219871 266085 219919 266113
rect 219609 266051 219919 266085
rect 219609 266023 219657 266051
rect 219685 266023 219719 266051
rect 219747 266023 219781 266051
rect 219809 266023 219843 266051
rect 219871 266023 219919 266051
rect 219609 265989 219919 266023
rect 219609 265961 219657 265989
rect 219685 265961 219719 265989
rect 219747 265961 219781 265989
rect 219809 265961 219843 265989
rect 219871 265961 219919 265989
rect 219609 257175 219919 265961
rect 219609 257147 219657 257175
rect 219685 257147 219719 257175
rect 219747 257147 219781 257175
rect 219809 257147 219843 257175
rect 219871 257147 219919 257175
rect 219609 257113 219919 257147
rect 219609 257085 219657 257113
rect 219685 257085 219719 257113
rect 219747 257085 219781 257113
rect 219809 257085 219843 257113
rect 219871 257085 219919 257113
rect 219609 257051 219919 257085
rect 219609 257023 219657 257051
rect 219685 257023 219719 257051
rect 219747 257023 219781 257051
rect 219809 257023 219843 257051
rect 219871 257023 219919 257051
rect 219609 256989 219919 257023
rect 219609 256961 219657 256989
rect 219685 256961 219719 256989
rect 219747 256961 219781 256989
rect 219809 256961 219843 256989
rect 219871 256961 219919 256989
rect 219609 248175 219919 256961
rect 219609 248147 219657 248175
rect 219685 248147 219719 248175
rect 219747 248147 219781 248175
rect 219809 248147 219843 248175
rect 219871 248147 219919 248175
rect 219609 248113 219919 248147
rect 219609 248085 219657 248113
rect 219685 248085 219719 248113
rect 219747 248085 219781 248113
rect 219809 248085 219843 248113
rect 219871 248085 219919 248113
rect 219609 248051 219919 248085
rect 219609 248023 219657 248051
rect 219685 248023 219719 248051
rect 219747 248023 219781 248051
rect 219809 248023 219843 248051
rect 219871 248023 219919 248051
rect 219609 247989 219919 248023
rect 219609 247961 219657 247989
rect 219685 247961 219719 247989
rect 219747 247961 219781 247989
rect 219809 247961 219843 247989
rect 219871 247961 219919 247989
rect 219609 239175 219919 247961
rect 219609 239147 219657 239175
rect 219685 239147 219719 239175
rect 219747 239147 219781 239175
rect 219809 239147 219843 239175
rect 219871 239147 219919 239175
rect 219609 239113 219919 239147
rect 219609 239085 219657 239113
rect 219685 239085 219719 239113
rect 219747 239085 219781 239113
rect 219809 239085 219843 239113
rect 219871 239085 219919 239113
rect 219609 239051 219919 239085
rect 219609 239023 219657 239051
rect 219685 239023 219719 239051
rect 219747 239023 219781 239051
rect 219809 239023 219843 239051
rect 219871 239023 219919 239051
rect 219609 238989 219919 239023
rect 219609 238961 219657 238989
rect 219685 238961 219719 238989
rect 219747 238961 219781 238989
rect 219809 238961 219843 238989
rect 219871 238961 219919 238989
rect 219609 230175 219919 238961
rect 219609 230147 219657 230175
rect 219685 230147 219719 230175
rect 219747 230147 219781 230175
rect 219809 230147 219843 230175
rect 219871 230147 219919 230175
rect 219609 230113 219919 230147
rect 219609 230085 219657 230113
rect 219685 230085 219719 230113
rect 219747 230085 219781 230113
rect 219809 230085 219843 230113
rect 219871 230085 219919 230113
rect 219609 230051 219919 230085
rect 219609 230023 219657 230051
rect 219685 230023 219719 230051
rect 219747 230023 219781 230051
rect 219809 230023 219843 230051
rect 219871 230023 219919 230051
rect 219609 229989 219919 230023
rect 219609 229961 219657 229989
rect 219685 229961 219719 229989
rect 219747 229961 219781 229989
rect 219809 229961 219843 229989
rect 219871 229961 219919 229989
rect 219609 221175 219919 229961
rect 219609 221147 219657 221175
rect 219685 221147 219719 221175
rect 219747 221147 219781 221175
rect 219809 221147 219843 221175
rect 219871 221147 219919 221175
rect 219609 221113 219919 221147
rect 219609 221085 219657 221113
rect 219685 221085 219719 221113
rect 219747 221085 219781 221113
rect 219809 221085 219843 221113
rect 219871 221085 219919 221113
rect 219609 221051 219919 221085
rect 219609 221023 219657 221051
rect 219685 221023 219719 221051
rect 219747 221023 219781 221051
rect 219809 221023 219843 221051
rect 219871 221023 219919 221051
rect 219609 220989 219919 221023
rect 219609 220961 219657 220989
rect 219685 220961 219719 220989
rect 219747 220961 219781 220989
rect 219809 220961 219843 220989
rect 219871 220961 219919 220989
rect 219609 212175 219919 220961
rect 219609 212147 219657 212175
rect 219685 212147 219719 212175
rect 219747 212147 219781 212175
rect 219809 212147 219843 212175
rect 219871 212147 219919 212175
rect 219609 212113 219919 212147
rect 219609 212085 219657 212113
rect 219685 212085 219719 212113
rect 219747 212085 219781 212113
rect 219809 212085 219843 212113
rect 219871 212085 219919 212113
rect 219609 212051 219919 212085
rect 219609 212023 219657 212051
rect 219685 212023 219719 212051
rect 219747 212023 219781 212051
rect 219809 212023 219843 212051
rect 219871 212023 219919 212051
rect 219609 211989 219919 212023
rect 219609 211961 219657 211989
rect 219685 211961 219719 211989
rect 219747 211961 219781 211989
rect 219809 211961 219843 211989
rect 219871 211961 219919 211989
rect 219609 203175 219919 211961
rect 219609 203147 219657 203175
rect 219685 203147 219719 203175
rect 219747 203147 219781 203175
rect 219809 203147 219843 203175
rect 219871 203147 219919 203175
rect 219609 203113 219919 203147
rect 219609 203085 219657 203113
rect 219685 203085 219719 203113
rect 219747 203085 219781 203113
rect 219809 203085 219843 203113
rect 219871 203085 219919 203113
rect 219609 203051 219919 203085
rect 219609 203023 219657 203051
rect 219685 203023 219719 203051
rect 219747 203023 219781 203051
rect 219809 203023 219843 203051
rect 219871 203023 219919 203051
rect 219609 202989 219919 203023
rect 219609 202961 219657 202989
rect 219685 202961 219719 202989
rect 219747 202961 219781 202989
rect 219809 202961 219843 202989
rect 219871 202961 219919 202989
rect 219609 194175 219919 202961
rect 219609 194147 219657 194175
rect 219685 194147 219719 194175
rect 219747 194147 219781 194175
rect 219809 194147 219843 194175
rect 219871 194147 219919 194175
rect 219609 194113 219919 194147
rect 219609 194085 219657 194113
rect 219685 194085 219719 194113
rect 219747 194085 219781 194113
rect 219809 194085 219843 194113
rect 219871 194085 219919 194113
rect 219609 194051 219919 194085
rect 219609 194023 219657 194051
rect 219685 194023 219719 194051
rect 219747 194023 219781 194051
rect 219809 194023 219843 194051
rect 219871 194023 219919 194051
rect 219609 193989 219919 194023
rect 219609 193961 219657 193989
rect 219685 193961 219719 193989
rect 219747 193961 219781 193989
rect 219809 193961 219843 193989
rect 219871 193961 219919 193989
rect 219609 185175 219919 193961
rect 219609 185147 219657 185175
rect 219685 185147 219719 185175
rect 219747 185147 219781 185175
rect 219809 185147 219843 185175
rect 219871 185147 219919 185175
rect 219609 185113 219919 185147
rect 219609 185085 219657 185113
rect 219685 185085 219719 185113
rect 219747 185085 219781 185113
rect 219809 185085 219843 185113
rect 219871 185085 219919 185113
rect 219609 185051 219919 185085
rect 219609 185023 219657 185051
rect 219685 185023 219719 185051
rect 219747 185023 219781 185051
rect 219809 185023 219843 185051
rect 219871 185023 219919 185051
rect 219609 184989 219919 185023
rect 219609 184961 219657 184989
rect 219685 184961 219719 184989
rect 219747 184961 219781 184989
rect 219809 184961 219843 184989
rect 219871 184961 219919 184989
rect 219609 176175 219919 184961
rect 219609 176147 219657 176175
rect 219685 176147 219719 176175
rect 219747 176147 219781 176175
rect 219809 176147 219843 176175
rect 219871 176147 219919 176175
rect 219609 176113 219919 176147
rect 219609 176085 219657 176113
rect 219685 176085 219719 176113
rect 219747 176085 219781 176113
rect 219809 176085 219843 176113
rect 219871 176085 219919 176113
rect 219609 176051 219919 176085
rect 219609 176023 219657 176051
rect 219685 176023 219719 176051
rect 219747 176023 219781 176051
rect 219809 176023 219843 176051
rect 219871 176023 219919 176051
rect 219609 175989 219919 176023
rect 219609 175961 219657 175989
rect 219685 175961 219719 175989
rect 219747 175961 219781 175989
rect 219809 175961 219843 175989
rect 219871 175961 219919 175989
rect 219609 167175 219919 175961
rect 219609 167147 219657 167175
rect 219685 167147 219719 167175
rect 219747 167147 219781 167175
rect 219809 167147 219843 167175
rect 219871 167147 219919 167175
rect 219609 167113 219919 167147
rect 219609 167085 219657 167113
rect 219685 167085 219719 167113
rect 219747 167085 219781 167113
rect 219809 167085 219843 167113
rect 219871 167085 219919 167113
rect 219609 167051 219919 167085
rect 219609 167023 219657 167051
rect 219685 167023 219719 167051
rect 219747 167023 219781 167051
rect 219809 167023 219843 167051
rect 219871 167023 219919 167051
rect 219609 166989 219919 167023
rect 219609 166961 219657 166989
rect 219685 166961 219719 166989
rect 219747 166961 219781 166989
rect 219809 166961 219843 166989
rect 219871 166961 219919 166989
rect 219609 158175 219919 166961
rect 233109 298606 233419 299134
rect 233109 298578 233157 298606
rect 233185 298578 233219 298606
rect 233247 298578 233281 298606
rect 233309 298578 233343 298606
rect 233371 298578 233419 298606
rect 233109 298544 233419 298578
rect 233109 298516 233157 298544
rect 233185 298516 233219 298544
rect 233247 298516 233281 298544
rect 233309 298516 233343 298544
rect 233371 298516 233419 298544
rect 233109 298482 233419 298516
rect 233109 298454 233157 298482
rect 233185 298454 233219 298482
rect 233247 298454 233281 298482
rect 233309 298454 233343 298482
rect 233371 298454 233419 298482
rect 233109 298420 233419 298454
rect 233109 298392 233157 298420
rect 233185 298392 233219 298420
rect 233247 298392 233281 298420
rect 233309 298392 233343 298420
rect 233371 298392 233419 298420
rect 233109 290175 233419 298392
rect 233109 290147 233157 290175
rect 233185 290147 233219 290175
rect 233247 290147 233281 290175
rect 233309 290147 233343 290175
rect 233371 290147 233419 290175
rect 233109 290113 233419 290147
rect 233109 290085 233157 290113
rect 233185 290085 233219 290113
rect 233247 290085 233281 290113
rect 233309 290085 233343 290113
rect 233371 290085 233419 290113
rect 233109 290051 233419 290085
rect 233109 290023 233157 290051
rect 233185 290023 233219 290051
rect 233247 290023 233281 290051
rect 233309 290023 233343 290051
rect 233371 290023 233419 290051
rect 233109 289989 233419 290023
rect 233109 289961 233157 289989
rect 233185 289961 233219 289989
rect 233247 289961 233281 289989
rect 233309 289961 233343 289989
rect 233371 289961 233419 289989
rect 233109 281175 233419 289961
rect 233109 281147 233157 281175
rect 233185 281147 233219 281175
rect 233247 281147 233281 281175
rect 233309 281147 233343 281175
rect 233371 281147 233419 281175
rect 233109 281113 233419 281147
rect 233109 281085 233157 281113
rect 233185 281085 233219 281113
rect 233247 281085 233281 281113
rect 233309 281085 233343 281113
rect 233371 281085 233419 281113
rect 233109 281051 233419 281085
rect 233109 281023 233157 281051
rect 233185 281023 233219 281051
rect 233247 281023 233281 281051
rect 233309 281023 233343 281051
rect 233371 281023 233419 281051
rect 233109 280989 233419 281023
rect 233109 280961 233157 280989
rect 233185 280961 233219 280989
rect 233247 280961 233281 280989
rect 233309 280961 233343 280989
rect 233371 280961 233419 280989
rect 233109 272175 233419 280961
rect 233109 272147 233157 272175
rect 233185 272147 233219 272175
rect 233247 272147 233281 272175
rect 233309 272147 233343 272175
rect 233371 272147 233419 272175
rect 233109 272113 233419 272147
rect 233109 272085 233157 272113
rect 233185 272085 233219 272113
rect 233247 272085 233281 272113
rect 233309 272085 233343 272113
rect 233371 272085 233419 272113
rect 233109 272051 233419 272085
rect 233109 272023 233157 272051
rect 233185 272023 233219 272051
rect 233247 272023 233281 272051
rect 233309 272023 233343 272051
rect 233371 272023 233419 272051
rect 233109 271989 233419 272023
rect 233109 271961 233157 271989
rect 233185 271961 233219 271989
rect 233247 271961 233281 271989
rect 233309 271961 233343 271989
rect 233371 271961 233419 271989
rect 233109 263175 233419 271961
rect 233109 263147 233157 263175
rect 233185 263147 233219 263175
rect 233247 263147 233281 263175
rect 233309 263147 233343 263175
rect 233371 263147 233419 263175
rect 233109 263113 233419 263147
rect 233109 263085 233157 263113
rect 233185 263085 233219 263113
rect 233247 263085 233281 263113
rect 233309 263085 233343 263113
rect 233371 263085 233419 263113
rect 233109 263051 233419 263085
rect 233109 263023 233157 263051
rect 233185 263023 233219 263051
rect 233247 263023 233281 263051
rect 233309 263023 233343 263051
rect 233371 263023 233419 263051
rect 233109 262989 233419 263023
rect 233109 262961 233157 262989
rect 233185 262961 233219 262989
rect 233247 262961 233281 262989
rect 233309 262961 233343 262989
rect 233371 262961 233419 262989
rect 233109 254175 233419 262961
rect 233109 254147 233157 254175
rect 233185 254147 233219 254175
rect 233247 254147 233281 254175
rect 233309 254147 233343 254175
rect 233371 254147 233419 254175
rect 233109 254113 233419 254147
rect 233109 254085 233157 254113
rect 233185 254085 233219 254113
rect 233247 254085 233281 254113
rect 233309 254085 233343 254113
rect 233371 254085 233419 254113
rect 233109 254051 233419 254085
rect 233109 254023 233157 254051
rect 233185 254023 233219 254051
rect 233247 254023 233281 254051
rect 233309 254023 233343 254051
rect 233371 254023 233419 254051
rect 233109 253989 233419 254023
rect 233109 253961 233157 253989
rect 233185 253961 233219 253989
rect 233247 253961 233281 253989
rect 233309 253961 233343 253989
rect 233371 253961 233419 253989
rect 233109 245175 233419 253961
rect 233109 245147 233157 245175
rect 233185 245147 233219 245175
rect 233247 245147 233281 245175
rect 233309 245147 233343 245175
rect 233371 245147 233419 245175
rect 233109 245113 233419 245147
rect 233109 245085 233157 245113
rect 233185 245085 233219 245113
rect 233247 245085 233281 245113
rect 233309 245085 233343 245113
rect 233371 245085 233419 245113
rect 233109 245051 233419 245085
rect 233109 245023 233157 245051
rect 233185 245023 233219 245051
rect 233247 245023 233281 245051
rect 233309 245023 233343 245051
rect 233371 245023 233419 245051
rect 233109 244989 233419 245023
rect 233109 244961 233157 244989
rect 233185 244961 233219 244989
rect 233247 244961 233281 244989
rect 233309 244961 233343 244989
rect 233371 244961 233419 244989
rect 233109 236175 233419 244961
rect 233109 236147 233157 236175
rect 233185 236147 233219 236175
rect 233247 236147 233281 236175
rect 233309 236147 233343 236175
rect 233371 236147 233419 236175
rect 233109 236113 233419 236147
rect 233109 236085 233157 236113
rect 233185 236085 233219 236113
rect 233247 236085 233281 236113
rect 233309 236085 233343 236113
rect 233371 236085 233419 236113
rect 233109 236051 233419 236085
rect 233109 236023 233157 236051
rect 233185 236023 233219 236051
rect 233247 236023 233281 236051
rect 233309 236023 233343 236051
rect 233371 236023 233419 236051
rect 233109 235989 233419 236023
rect 233109 235961 233157 235989
rect 233185 235961 233219 235989
rect 233247 235961 233281 235989
rect 233309 235961 233343 235989
rect 233371 235961 233419 235989
rect 233109 227175 233419 235961
rect 233109 227147 233157 227175
rect 233185 227147 233219 227175
rect 233247 227147 233281 227175
rect 233309 227147 233343 227175
rect 233371 227147 233419 227175
rect 233109 227113 233419 227147
rect 233109 227085 233157 227113
rect 233185 227085 233219 227113
rect 233247 227085 233281 227113
rect 233309 227085 233343 227113
rect 233371 227085 233419 227113
rect 233109 227051 233419 227085
rect 233109 227023 233157 227051
rect 233185 227023 233219 227051
rect 233247 227023 233281 227051
rect 233309 227023 233343 227051
rect 233371 227023 233419 227051
rect 233109 226989 233419 227023
rect 233109 226961 233157 226989
rect 233185 226961 233219 226989
rect 233247 226961 233281 226989
rect 233309 226961 233343 226989
rect 233371 226961 233419 226989
rect 233109 218175 233419 226961
rect 233109 218147 233157 218175
rect 233185 218147 233219 218175
rect 233247 218147 233281 218175
rect 233309 218147 233343 218175
rect 233371 218147 233419 218175
rect 233109 218113 233419 218147
rect 233109 218085 233157 218113
rect 233185 218085 233219 218113
rect 233247 218085 233281 218113
rect 233309 218085 233343 218113
rect 233371 218085 233419 218113
rect 233109 218051 233419 218085
rect 233109 218023 233157 218051
rect 233185 218023 233219 218051
rect 233247 218023 233281 218051
rect 233309 218023 233343 218051
rect 233371 218023 233419 218051
rect 233109 217989 233419 218023
rect 233109 217961 233157 217989
rect 233185 217961 233219 217989
rect 233247 217961 233281 217989
rect 233309 217961 233343 217989
rect 233371 217961 233419 217989
rect 233109 209175 233419 217961
rect 233109 209147 233157 209175
rect 233185 209147 233219 209175
rect 233247 209147 233281 209175
rect 233309 209147 233343 209175
rect 233371 209147 233419 209175
rect 233109 209113 233419 209147
rect 233109 209085 233157 209113
rect 233185 209085 233219 209113
rect 233247 209085 233281 209113
rect 233309 209085 233343 209113
rect 233371 209085 233419 209113
rect 233109 209051 233419 209085
rect 233109 209023 233157 209051
rect 233185 209023 233219 209051
rect 233247 209023 233281 209051
rect 233309 209023 233343 209051
rect 233371 209023 233419 209051
rect 233109 208989 233419 209023
rect 233109 208961 233157 208989
rect 233185 208961 233219 208989
rect 233247 208961 233281 208989
rect 233309 208961 233343 208989
rect 233371 208961 233419 208989
rect 233109 200175 233419 208961
rect 233109 200147 233157 200175
rect 233185 200147 233219 200175
rect 233247 200147 233281 200175
rect 233309 200147 233343 200175
rect 233371 200147 233419 200175
rect 233109 200113 233419 200147
rect 233109 200085 233157 200113
rect 233185 200085 233219 200113
rect 233247 200085 233281 200113
rect 233309 200085 233343 200113
rect 233371 200085 233419 200113
rect 233109 200051 233419 200085
rect 233109 200023 233157 200051
rect 233185 200023 233219 200051
rect 233247 200023 233281 200051
rect 233309 200023 233343 200051
rect 233371 200023 233419 200051
rect 233109 199989 233419 200023
rect 233109 199961 233157 199989
rect 233185 199961 233219 199989
rect 233247 199961 233281 199989
rect 233309 199961 233343 199989
rect 233371 199961 233419 199989
rect 233109 191175 233419 199961
rect 233109 191147 233157 191175
rect 233185 191147 233219 191175
rect 233247 191147 233281 191175
rect 233309 191147 233343 191175
rect 233371 191147 233419 191175
rect 233109 191113 233419 191147
rect 233109 191085 233157 191113
rect 233185 191085 233219 191113
rect 233247 191085 233281 191113
rect 233309 191085 233343 191113
rect 233371 191085 233419 191113
rect 233109 191051 233419 191085
rect 233109 191023 233157 191051
rect 233185 191023 233219 191051
rect 233247 191023 233281 191051
rect 233309 191023 233343 191051
rect 233371 191023 233419 191051
rect 233109 190989 233419 191023
rect 233109 190961 233157 190989
rect 233185 190961 233219 190989
rect 233247 190961 233281 190989
rect 233309 190961 233343 190989
rect 233371 190961 233419 190989
rect 233109 182175 233419 190961
rect 233109 182147 233157 182175
rect 233185 182147 233219 182175
rect 233247 182147 233281 182175
rect 233309 182147 233343 182175
rect 233371 182147 233419 182175
rect 233109 182113 233419 182147
rect 233109 182085 233157 182113
rect 233185 182085 233219 182113
rect 233247 182085 233281 182113
rect 233309 182085 233343 182113
rect 233371 182085 233419 182113
rect 233109 182051 233419 182085
rect 233109 182023 233157 182051
rect 233185 182023 233219 182051
rect 233247 182023 233281 182051
rect 233309 182023 233343 182051
rect 233371 182023 233419 182051
rect 233109 181989 233419 182023
rect 233109 181961 233157 181989
rect 233185 181961 233219 181989
rect 233247 181961 233281 181989
rect 233309 181961 233343 181989
rect 233371 181961 233419 181989
rect 233109 173175 233419 181961
rect 233109 173147 233157 173175
rect 233185 173147 233219 173175
rect 233247 173147 233281 173175
rect 233309 173147 233343 173175
rect 233371 173147 233419 173175
rect 233109 173113 233419 173147
rect 233109 173085 233157 173113
rect 233185 173085 233219 173113
rect 233247 173085 233281 173113
rect 233309 173085 233343 173113
rect 233371 173085 233419 173113
rect 233109 173051 233419 173085
rect 233109 173023 233157 173051
rect 233185 173023 233219 173051
rect 233247 173023 233281 173051
rect 233309 173023 233343 173051
rect 233371 173023 233419 173051
rect 233109 172989 233419 173023
rect 233109 172961 233157 172989
rect 233185 172961 233219 172989
rect 233247 172961 233281 172989
rect 233309 172961 233343 172989
rect 233371 172961 233419 172989
rect 233109 164175 233419 172961
rect 233109 164147 233157 164175
rect 233185 164147 233219 164175
rect 233247 164147 233281 164175
rect 233309 164147 233343 164175
rect 233371 164147 233419 164175
rect 233109 164113 233419 164147
rect 233109 164085 233157 164113
rect 233185 164085 233219 164113
rect 233247 164085 233281 164113
rect 233309 164085 233343 164113
rect 233371 164085 233419 164113
rect 233109 164051 233419 164085
rect 233109 164023 233157 164051
rect 233185 164023 233219 164051
rect 233247 164023 233281 164051
rect 233309 164023 233343 164051
rect 233371 164023 233419 164051
rect 233109 163989 233419 164023
rect 233109 163961 233157 163989
rect 233185 163961 233219 163989
rect 233247 163961 233281 163989
rect 233309 163961 233343 163989
rect 233371 163961 233419 163989
rect 219609 158147 219657 158175
rect 219685 158147 219719 158175
rect 219747 158147 219781 158175
rect 219809 158147 219843 158175
rect 219871 158147 219919 158175
rect 219609 158113 219919 158147
rect 219609 158085 219657 158113
rect 219685 158085 219719 158113
rect 219747 158085 219781 158113
rect 219809 158085 219843 158113
rect 219871 158085 219919 158113
rect 219609 158051 219919 158085
rect 219609 158023 219657 158051
rect 219685 158023 219719 158051
rect 219747 158023 219781 158051
rect 219809 158023 219843 158051
rect 219871 158023 219919 158051
rect 219609 157989 219919 158023
rect 219609 157961 219657 157989
rect 219685 157961 219719 157989
rect 219747 157961 219781 157989
rect 219809 157961 219843 157989
rect 219871 157961 219919 157989
rect 219609 149175 219919 157961
rect 224224 158175 224384 158192
rect 224224 158147 224259 158175
rect 224287 158147 224321 158175
rect 224349 158147 224384 158175
rect 224224 158113 224384 158147
rect 224224 158085 224259 158113
rect 224287 158085 224321 158113
rect 224349 158085 224384 158113
rect 224224 158051 224384 158085
rect 224224 158023 224259 158051
rect 224287 158023 224321 158051
rect 224349 158023 224384 158051
rect 224224 157989 224384 158023
rect 224224 157961 224259 157989
rect 224287 157961 224321 157989
rect 224349 157961 224384 157989
rect 224224 157944 224384 157961
rect 231904 155175 232064 155192
rect 231904 155147 231939 155175
rect 231967 155147 232001 155175
rect 232029 155147 232064 155175
rect 231904 155113 232064 155147
rect 231904 155085 231939 155113
rect 231967 155085 232001 155113
rect 232029 155085 232064 155113
rect 231904 155051 232064 155085
rect 231904 155023 231939 155051
rect 231967 155023 232001 155051
rect 232029 155023 232064 155051
rect 231904 154989 232064 155023
rect 231904 154961 231939 154989
rect 231967 154961 232001 154989
rect 232029 154961 232064 154989
rect 231904 154944 232064 154961
rect 233109 155175 233419 163961
rect 233109 155147 233157 155175
rect 233185 155147 233219 155175
rect 233247 155147 233281 155175
rect 233309 155147 233343 155175
rect 233371 155147 233419 155175
rect 233109 155113 233419 155147
rect 233109 155085 233157 155113
rect 233185 155085 233219 155113
rect 233247 155085 233281 155113
rect 233309 155085 233343 155113
rect 233371 155085 233419 155113
rect 233109 155051 233419 155085
rect 233109 155023 233157 155051
rect 233185 155023 233219 155051
rect 233247 155023 233281 155051
rect 233309 155023 233343 155051
rect 233371 155023 233419 155051
rect 233109 154989 233419 155023
rect 233109 154961 233157 154989
rect 233185 154961 233219 154989
rect 233247 154961 233281 154989
rect 233309 154961 233343 154989
rect 233371 154961 233419 154989
rect 219609 149147 219657 149175
rect 219685 149147 219719 149175
rect 219747 149147 219781 149175
rect 219809 149147 219843 149175
rect 219871 149147 219919 149175
rect 219609 149113 219919 149147
rect 219609 149085 219657 149113
rect 219685 149085 219719 149113
rect 219747 149085 219781 149113
rect 219809 149085 219843 149113
rect 219871 149085 219919 149113
rect 219609 149051 219919 149085
rect 219609 149023 219657 149051
rect 219685 149023 219719 149051
rect 219747 149023 219781 149051
rect 219809 149023 219843 149051
rect 219871 149023 219919 149051
rect 219609 148989 219919 149023
rect 219609 148961 219657 148989
rect 219685 148961 219719 148989
rect 219747 148961 219781 148989
rect 219809 148961 219843 148989
rect 219871 148961 219919 148989
rect 219609 140175 219919 148961
rect 224224 149175 224384 149192
rect 224224 149147 224259 149175
rect 224287 149147 224321 149175
rect 224349 149147 224384 149175
rect 224224 149113 224384 149147
rect 224224 149085 224259 149113
rect 224287 149085 224321 149113
rect 224349 149085 224384 149113
rect 224224 149051 224384 149085
rect 224224 149023 224259 149051
rect 224287 149023 224321 149051
rect 224349 149023 224384 149051
rect 224224 148989 224384 149023
rect 224224 148961 224259 148989
rect 224287 148961 224321 148989
rect 224349 148961 224384 148989
rect 224224 148944 224384 148961
rect 231904 146175 232064 146192
rect 231904 146147 231939 146175
rect 231967 146147 232001 146175
rect 232029 146147 232064 146175
rect 231904 146113 232064 146147
rect 231904 146085 231939 146113
rect 231967 146085 232001 146113
rect 232029 146085 232064 146113
rect 231904 146051 232064 146085
rect 231904 146023 231939 146051
rect 231967 146023 232001 146051
rect 232029 146023 232064 146051
rect 231904 145989 232064 146023
rect 231904 145961 231939 145989
rect 231967 145961 232001 145989
rect 232029 145961 232064 145989
rect 231904 145944 232064 145961
rect 233109 146175 233419 154961
rect 233109 146147 233157 146175
rect 233185 146147 233219 146175
rect 233247 146147 233281 146175
rect 233309 146147 233343 146175
rect 233371 146147 233419 146175
rect 233109 146113 233419 146147
rect 233109 146085 233157 146113
rect 233185 146085 233219 146113
rect 233247 146085 233281 146113
rect 233309 146085 233343 146113
rect 233371 146085 233419 146113
rect 233109 146051 233419 146085
rect 233109 146023 233157 146051
rect 233185 146023 233219 146051
rect 233247 146023 233281 146051
rect 233309 146023 233343 146051
rect 233371 146023 233419 146051
rect 233109 145989 233419 146023
rect 233109 145961 233157 145989
rect 233185 145961 233219 145989
rect 233247 145961 233281 145989
rect 233309 145961 233343 145989
rect 233371 145961 233419 145989
rect 219609 140147 219657 140175
rect 219685 140147 219719 140175
rect 219747 140147 219781 140175
rect 219809 140147 219843 140175
rect 219871 140147 219919 140175
rect 219609 140113 219919 140147
rect 219609 140085 219657 140113
rect 219685 140085 219719 140113
rect 219747 140085 219781 140113
rect 219809 140085 219843 140113
rect 219871 140085 219919 140113
rect 219609 140051 219919 140085
rect 219609 140023 219657 140051
rect 219685 140023 219719 140051
rect 219747 140023 219781 140051
rect 219809 140023 219843 140051
rect 219871 140023 219919 140051
rect 219609 139989 219919 140023
rect 219609 139961 219657 139989
rect 219685 139961 219719 139989
rect 219747 139961 219781 139989
rect 219809 139961 219843 139989
rect 219871 139961 219919 139989
rect 219609 131175 219919 139961
rect 224224 140175 224384 140192
rect 224224 140147 224259 140175
rect 224287 140147 224321 140175
rect 224349 140147 224384 140175
rect 224224 140113 224384 140147
rect 224224 140085 224259 140113
rect 224287 140085 224321 140113
rect 224349 140085 224384 140113
rect 224224 140051 224384 140085
rect 224224 140023 224259 140051
rect 224287 140023 224321 140051
rect 224349 140023 224384 140051
rect 224224 139989 224384 140023
rect 224224 139961 224259 139989
rect 224287 139961 224321 139989
rect 224349 139961 224384 139989
rect 224224 139944 224384 139961
rect 231904 137175 232064 137192
rect 231904 137147 231939 137175
rect 231967 137147 232001 137175
rect 232029 137147 232064 137175
rect 231904 137113 232064 137147
rect 231904 137085 231939 137113
rect 231967 137085 232001 137113
rect 232029 137085 232064 137113
rect 231904 137051 232064 137085
rect 231904 137023 231939 137051
rect 231967 137023 232001 137051
rect 232029 137023 232064 137051
rect 231904 136989 232064 137023
rect 231904 136961 231939 136989
rect 231967 136961 232001 136989
rect 232029 136961 232064 136989
rect 231904 136944 232064 136961
rect 233109 137175 233419 145961
rect 233109 137147 233157 137175
rect 233185 137147 233219 137175
rect 233247 137147 233281 137175
rect 233309 137147 233343 137175
rect 233371 137147 233419 137175
rect 233109 137113 233419 137147
rect 233109 137085 233157 137113
rect 233185 137085 233219 137113
rect 233247 137085 233281 137113
rect 233309 137085 233343 137113
rect 233371 137085 233419 137113
rect 233109 137051 233419 137085
rect 233109 137023 233157 137051
rect 233185 137023 233219 137051
rect 233247 137023 233281 137051
rect 233309 137023 233343 137051
rect 233371 137023 233419 137051
rect 233109 136989 233419 137023
rect 233109 136961 233157 136989
rect 233185 136961 233219 136989
rect 233247 136961 233281 136989
rect 233309 136961 233343 136989
rect 233371 136961 233419 136989
rect 219609 131147 219657 131175
rect 219685 131147 219719 131175
rect 219747 131147 219781 131175
rect 219809 131147 219843 131175
rect 219871 131147 219919 131175
rect 219609 131113 219919 131147
rect 219609 131085 219657 131113
rect 219685 131085 219719 131113
rect 219747 131085 219781 131113
rect 219809 131085 219843 131113
rect 219871 131085 219919 131113
rect 219609 131051 219919 131085
rect 219609 131023 219657 131051
rect 219685 131023 219719 131051
rect 219747 131023 219781 131051
rect 219809 131023 219843 131051
rect 219871 131023 219919 131051
rect 219609 130989 219919 131023
rect 219609 130961 219657 130989
rect 219685 130961 219719 130989
rect 219747 130961 219781 130989
rect 219809 130961 219843 130989
rect 219871 130961 219919 130989
rect 219609 125367 219919 130961
rect 233109 128175 233419 136961
rect 233109 128147 233157 128175
rect 233185 128147 233219 128175
rect 233247 128147 233281 128175
rect 233309 128147 233343 128175
rect 233371 128147 233419 128175
rect 233109 128113 233419 128147
rect 233109 128085 233157 128113
rect 233185 128085 233219 128113
rect 233247 128085 233281 128113
rect 233309 128085 233343 128113
rect 233371 128085 233419 128113
rect 233109 128051 233419 128085
rect 233109 128023 233157 128051
rect 233185 128023 233219 128051
rect 233247 128023 233281 128051
rect 233309 128023 233343 128051
rect 233371 128023 233419 128051
rect 233109 127989 233419 128023
rect 233109 127961 233157 127989
rect 233185 127961 233219 127989
rect 233247 127961 233281 127989
rect 233309 127961 233343 127989
rect 233371 127961 233419 127989
rect 233109 125367 233419 127961
rect 234969 299086 235279 299134
rect 234969 299058 235017 299086
rect 235045 299058 235079 299086
rect 235107 299058 235141 299086
rect 235169 299058 235203 299086
rect 235231 299058 235279 299086
rect 234969 299024 235279 299058
rect 234969 298996 235017 299024
rect 235045 298996 235079 299024
rect 235107 298996 235141 299024
rect 235169 298996 235203 299024
rect 235231 298996 235279 299024
rect 234969 298962 235279 298996
rect 234969 298934 235017 298962
rect 235045 298934 235079 298962
rect 235107 298934 235141 298962
rect 235169 298934 235203 298962
rect 235231 298934 235279 298962
rect 234969 298900 235279 298934
rect 234969 298872 235017 298900
rect 235045 298872 235079 298900
rect 235107 298872 235141 298900
rect 235169 298872 235203 298900
rect 235231 298872 235279 298900
rect 234969 293175 235279 298872
rect 234969 293147 235017 293175
rect 235045 293147 235079 293175
rect 235107 293147 235141 293175
rect 235169 293147 235203 293175
rect 235231 293147 235279 293175
rect 234969 293113 235279 293147
rect 234969 293085 235017 293113
rect 235045 293085 235079 293113
rect 235107 293085 235141 293113
rect 235169 293085 235203 293113
rect 235231 293085 235279 293113
rect 234969 293051 235279 293085
rect 234969 293023 235017 293051
rect 235045 293023 235079 293051
rect 235107 293023 235141 293051
rect 235169 293023 235203 293051
rect 235231 293023 235279 293051
rect 234969 292989 235279 293023
rect 234969 292961 235017 292989
rect 235045 292961 235079 292989
rect 235107 292961 235141 292989
rect 235169 292961 235203 292989
rect 235231 292961 235279 292989
rect 234969 284175 235279 292961
rect 234969 284147 235017 284175
rect 235045 284147 235079 284175
rect 235107 284147 235141 284175
rect 235169 284147 235203 284175
rect 235231 284147 235279 284175
rect 234969 284113 235279 284147
rect 234969 284085 235017 284113
rect 235045 284085 235079 284113
rect 235107 284085 235141 284113
rect 235169 284085 235203 284113
rect 235231 284085 235279 284113
rect 234969 284051 235279 284085
rect 234969 284023 235017 284051
rect 235045 284023 235079 284051
rect 235107 284023 235141 284051
rect 235169 284023 235203 284051
rect 235231 284023 235279 284051
rect 234969 283989 235279 284023
rect 234969 283961 235017 283989
rect 235045 283961 235079 283989
rect 235107 283961 235141 283989
rect 235169 283961 235203 283989
rect 235231 283961 235279 283989
rect 234969 275175 235279 283961
rect 234969 275147 235017 275175
rect 235045 275147 235079 275175
rect 235107 275147 235141 275175
rect 235169 275147 235203 275175
rect 235231 275147 235279 275175
rect 234969 275113 235279 275147
rect 234969 275085 235017 275113
rect 235045 275085 235079 275113
rect 235107 275085 235141 275113
rect 235169 275085 235203 275113
rect 235231 275085 235279 275113
rect 234969 275051 235279 275085
rect 234969 275023 235017 275051
rect 235045 275023 235079 275051
rect 235107 275023 235141 275051
rect 235169 275023 235203 275051
rect 235231 275023 235279 275051
rect 234969 274989 235279 275023
rect 234969 274961 235017 274989
rect 235045 274961 235079 274989
rect 235107 274961 235141 274989
rect 235169 274961 235203 274989
rect 235231 274961 235279 274989
rect 234969 266175 235279 274961
rect 234969 266147 235017 266175
rect 235045 266147 235079 266175
rect 235107 266147 235141 266175
rect 235169 266147 235203 266175
rect 235231 266147 235279 266175
rect 234969 266113 235279 266147
rect 234969 266085 235017 266113
rect 235045 266085 235079 266113
rect 235107 266085 235141 266113
rect 235169 266085 235203 266113
rect 235231 266085 235279 266113
rect 234969 266051 235279 266085
rect 234969 266023 235017 266051
rect 235045 266023 235079 266051
rect 235107 266023 235141 266051
rect 235169 266023 235203 266051
rect 235231 266023 235279 266051
rect 234969 265989 235279 266023
rect 234969 265961 235017 265989
rect 235045 265961 235079 265989
rect 235107 265961 235141 265989
rect 235169 265961 235203 265989
rect 235231 265961 235279 265989
rect 234969 257175 235279 265961
rect 234969 257147 235017 257175
rect 235045 257147 235079 257175
rect 235107 257147 235141 257175
rect 235169 257147 235203 257175
rect 235231 257147 235279 257175
rect 234969 257113 235279 257147
rect 234969 257085 235017 257113
rect 235045 257085 235079 257113
rect 235107 257085 235141 257113
rect 235169 257085 235203 257113
rect 235231 257085 235279 257113
rect 234969 257051 235279 257085
rect 234969 257023 235017 257051
rect 235045 257023 235079 257051
rect 235107 257023 235141 257051
rect 235169 257023 235203 257051
rect 235231 257023 235279 257051
rect 234969 256989 235279 257023
rect 234969 256961 235017 256989
rect 235045 256961 235079 256989
rect 235107 256961 235141 256989
rect 235169 256961 235203 256989
rect 235231 256961 235279 256989
rect 234969 248175 235279 256961
rect 234969 248147 235017 248175
rect 235045 248147 235079 248175
rect 235107 248147 235141 248175
rect 235169 248147 235203 248175
rect 235231 248147 235279 248175
rect 234969 248113 235279 248147
rect 234969 248085 235017 248113
rect 235045 248085 235079 248113
rect 235107 248085 235141 248113
rect 235169 248085 235203 248113
rect 235231 248085 235279 248113
rect 234969 248051 235279 248085
rect 234969 248023 235017 248051
rect 235045 248023 235079 248051
rect 235107 248023 235141 248051
rect 235169 248023 235203 248051
rect 235231 248023 235279 248051
rect 234969 247989 235279 248023
rect 234969 247961 235017 247989
rect 235045 247961 235079 247989
rect 235107 247961 235141 247989
rect 235169 247961 235203 247989
rect 235231 247961 235279 247989
rect 234969 239175 235279 247961
rect 234969 239147 235017 239175
rect 235045 239147 235079 239175
rect 235107 239147 235141 239175
rect 235169 239147 235203 239175
rect 235231 239147 235279 239175
rect 234969 239113 235279 239147
rect 234969 239085 235017 239113
rect 235045 239085 235079 239113
rect 235107 239085 235141 239113
rect 235169 239085 235203 239113
rect 235231 239085 235279 239113
rect 234969 239051 235279 239085
rect 234969 239023 235017 239051
rect 235045 239023 235079 239051
rect 235107 239023 235141 239051
rect 235169 239023 235203 239051
rect 235231 239023 235279 239051
rect 234969 238989 235279 239023
rect 234969 238961 235017 238989
rect 235045 238961 235079 238989
rect 235107 238961 235141 238989
rect 235169 238961 235203 238989
rect 235231 238961 235279 238989
rect 234969 230175 235279 238961
rect 234969 230147 235017 230175
rect 235045 230147 235079 230175
rect 235107 230147 235141 230175
rect 235169 230147 235203 230175
rect 235231 230147 235279 230175
rect 234969 230113 235279 230147
rect 234969 230085 235017 230113
rect 235045 230085 235079 230113
rect 235107 230085 235141 230113
rect 235169 230085 235203 230113
rect 235231 230085 235279 230113
rect 234969 230051 235279 230085
rect 234969 230023 235017 230051
rect 235045 230023 235079 230051
rect 235107 230023 235141 230051
rect 235169 230023 235203 230051
rect 235231 230023 235279 230051
rect 234969 229989 235279 230023
rect 234969 229961 235017 229989
rect 235045 229961 235079 229989
rect 235107 229961 235141 229989
rect 235169 229961 235203 229989
rect 235231 229961 235279 229989
rect 234969 221175 235279 229961
rect 234969 221147 235017 221175
rect 235045 221147 235079 221175
rect 235107 221147 235141 221175
rect 235169 221147 235203 221175
rect 235231 221147 235279 221175
rect 234969 221113 235279 221147
rect 234969 221085 235017 221113
rect 235045 221085 235079 221113
rect 235107 221085 235141 221113
rect 235169 221085 235203 221113
rect 235231 221085 235279 221113
rect 234969 221051 235279 221085
rect 234969 221023 235017 221051
rect 235045 221023 235079 221051
rect 235107 221023 235141 221051
rect 235169 221023 235203 221051
rect 235231 221023 235279 221051
rect 234969 220989 235279 221023
rect 234969 220961 235017 220989
rect 235045 220961 235079 220989
rect 235107 220961 235141 220989
rect 235169 220961 235203 220989
rect 235231 220961 235279 220989
rect 234969 212175 235279 220961
rect 234969 212147 235017 212175
rect 235045 212147 235079 212175
rect 235107 212147 235141 212175
rect 235169 212147 235203 212175
rect 235231 212147 235279 212175
rect 234969 212113 235279 212147
rect 234969 212085 235017 212113
rect 235045 212085 235079 212113
rect 235107 212085 235141 212113
rect 235169 212085 235203 212113
rect 235231 212085 235279 212113
rect 234969 212051 235279 212085
rect 234969 212023 235017 212051
rect 235045 212023 235079 212051
rect 235107 212023 235141 212051
rect 235169 212023 235203 212051
rect 235231 212023 235279 212051
rect 234969 211989 235279 212023
rect 234969 211961 235017 211989
rect 235045 211961 235079 211989
rect 235107 211961 235141 211989
rect 235169 211961 235203 211989
rect 235231 211961 235279 211989
rect 234969 203175 235279 211961
rect 234969 203147 235017 203175
rect 235045 203147 235079 203175
rect 235107 203147 235141 203175
rect 235169 203147 235203 203175
rect 235231 203147 235279 203175
rect 234969 203113 235279 203147
rect 234969 203085 235017 203113
rect 235045 203085 235079 203113
rect 235107 203085 235141 203113
rect 235169 203085 235203 203113
rect 235231 203085 235279 203113
rect 234969 203051 235279 203085
rect 234969 203023 235017 203051
rect 235045 203023 235079 203051
rect 235107 203023 235141 203051
rect 235169 203023 235203 203051
rect 235231 203023 235279 203051
rect 234969 202989 235279 203023
rect 234969 202961 235017 202989
rect 235045 202961 235079 202989
rect 235107 202961 235141 202989
rect 235169 202961 235203 202989
rect 235231 202961 235279 202989
rect 234969 194175 235279 202961
rect 234969 194147 235017 194175
rect 235045 194147 235079 194175
rect 235107 194147 235141 194175
rect 235169 194147 235203 194175
rect 235231 194147 235279 194175
rect 234969 194113 235279 194147
rect 234969 194085 235017 194113
rect 235045 194085 235079 194113
rect 235107 194085 235141 194113
rect 235169 194085 235203 194113
rect 235231 194085 235279 194113
rect 234969 194051 235279 194085
rect 234969 194023 235017 194051
rect 235045 194023 235079 194051
rect 235107 194023 235141 194051
rect 235169 194023 235203 194051
rect 235231 194023 235279 194051
rect 234969 193989 235279 194023
rect 234969 193961 235017 193989
rect 235045 193961 235079 193989
rect 235107 193961 235141 193989
rect 235169 193961 235203 193989
rect 235231 193961 235279 193989
rect 234969 185175 235279 193961
rect 248469 298606 248779 299134
rect 248469 298578 248517 298606
rect 248545 298578 248579 298606
rect 248607 298578 248641 298606
rect 248669 298578 248703 298606
rect 248731 298578 248779 298606
rect 248469 298544 248779 298578
rect 248469 298516 248517 298544
rect 248545 298516 248579 298544
rect 248607 298516 248641 298544
rect 248669 298516 248703 298544
rect 248731 298516 248779 298544
rect 248469 298482 248779 298516
rect 248469 298454 248517 298482
rect 248545 298454 248579 298482
rect 248607 298454 248641 298482
rect 248669 298454 248703 298482
rect 248731 298454 248779 298482
rect 248469 298420 248779 298454
rect 248469 298392 248517 298420
rect 248545 298392 248579 298420
rect 248607 298392 248641 298420
rect 248669 298392 248703 298420
rect 248731 298392 248779 298420
rect 248469 290175 248779 298392
rect 248469 290147 248517 290175
rect 248545 290147 248579 290175
rect 248607 290147 248641 290175
rect 248669 290147 248703 290175
rect 248731 290147 248779 290175
rect 248469 290113 248779 290147
rect 248469 290085 248517 290113
rect 248545 290085 248579 290113
rect 248607 290085 248641 290113
rect 248669 290085 248703 290113
rect 248731 290085 248779 290113
rect 248469 290051 248779 290085
rect 248469 290023 248517 290051
rect 248545 290023 248579 290051
rect 248607 290023 248641 290051
rect 248669 290023 248703 290051
rect 248731 290023 248779 290051
rect 248469 289989 248779 290023
rect 248469 289961 248517 289989
rect 248545 289961 248579 289989
rect 248607 289961 248641 289989
rect 248669 289961 248703 289989
rect 248731 289961 248779 289989
rect 248469 281175 248779 289961
rect 248469 281147 248517 281175
rect 248545 281147 248579 281175
rect 248607 281147 248641 281175
rect 248669 281147 248703 281175
rect 248731 281147 248779 281175
rect 248469 281113 248779 281147
rect 248469 281085 248517 281113
rect 248545 281085 248579 281113
rect 248607 281085 248641 281113
rect 248669 281085 248703 281113
rect 248731 281085 248779 281113
rect 248469 281051 248779 281085
rect 248469 281023 248517 281051
rect 248545 281023 248579 281051
rect 248607 281023 248641 281051
rect 248669 281023 248703 281051
rect 248731 281023 248779 281051
rect 248469 280989 248779 281023
rect 248469 280961 248517 280989
rect 248545 280961 248579 280989
rect 248607 280961 248641 280989
rect 248669 280961 248703 280989
rect 248731 280961 248779 280989
rect 248469 272175 248779 280961
rect 248469 272147 248517 272175
rect 248545 272147 248579 272175
rect 248607 272147 248641 272175
rect 248669 272147 248703 272175
rect 248731 272147 248779 272175
rect 248469 272113 248779 272147
rect 248469 272085 248517 272113
rect 248545 272085 248579 272113
rect 248607 272085 248641 272113
rect 248669 272085 248703 272113
rect 248731 272085 248779 272113
rect 248469 272051 248779 272085
rect 248469 272023 248517 272051
rect 248545 272023 248579 272051
rect 248607 272023 248641 272051
rect 248669 272023 248703 272051
rect 248731 272023 248779 272051
rect 248469 271989 248779 272023
rect 248469 271961 248517 271989
rect 248545 271961 248579 271989
rect 248607 271961 248641 271989
rect 248669 271961 248703 271989
rect 248731 271961 248779 271989
rect 248469 263175 248779 271961
rect 248469 263147 248517 263175
rect 248545 263147 248579 263175
rect 248607 263147 248641 263175
rect 248669 263147 248703 263175
rect 248731 263147 248779 263175
rect 248469 263113 248779 263147
rect 248469 263085 248517 263113
rect 248545 263085 248579 263113
rect 248607 263085 248641 263113
rect 248669 263085 248703 263113
rect 248731 263085 248779 263113
rect 248469 263051 248779 263085
rect 248469 263023 248517 263051
rect 248545 263023 248579 263051
rect 248607 263023 248641 263051
rect 248669 263023 248703 263051
rect 248731 263023 248779 263051
rect 248469 262989 248779 263023
rect 248469 262961 248517 262989
rect 248545 262961 248579 262989
rect 248607 262961 248641 262989
rect 248669 262961 248703 262989
rect 248731 262961 248779 262989
rect 248469 254175 248779 262961
rect 248469 254147 248517 254175
rect 248545 254147 248579 254175
rect 248607 254147 248641 254175
rect 248669 254147 248703 254175
rect 248731 254147 248779 254175
rect 248469 254113 248779 254147
rect 248469 254085 248517 254113
rect 248545 254085 248579 254113
rect 248607 254085 248641 254113
rect 248669 254085 248703 254113
rect 248731 254085 248779 254113
rect 248469 254051 248779 254085
rect 248469 254023 248517 254051
rect 248545 254023 248579 254051
rect 248607 254023 248641 254051
rect 248669 254023 248703 254051
rect 248731 254023 248779 254051
rect 248469 253989 248779 254023
rect 248469 253961 248517 253989
rect 248545 253961 248579 253989
rect 248607 253961 248641 253989
rect 248669 253961 248703 253989
rect 248731 253961 248779 253989
rect 248469 245175 248779 253961
rect 248469 245147 248517 245175
rect 248545 245147 248579 245175
rect 248607 245147 248641 245175
rect 248669 245147 248703 245175
rect 248731 245147 248779 245175
rect 248469 245113 248779 245147
rect 248469 245085 248517 245113
rect 248545 245085 248579 245113
rect 248607 245085 248641 245113
rect 248669 245085 248703 245113
rect 248731 245085 248779 245113
rect 248469 245051 248779 245085
rect 248469 245023 248517 245051
rect 248545 245023 248579 245051
rect 248607 245023 248641 245051
rect 248669 245023 248703 245051
rect 248731 245023 248779 245051
rect 248469 244989 248779 245023
rect 248469 244961 248517 244989
rect 248545 244961 248579 244989
rect 248607 244961 248641 244989
rect 248669 244961 248703 244989
rect 248731 244961 248779 244989
rect 248469 236175 248779 244961
rect 248469 236147 248517 236175
rect 248545 236147 248579 236175
rect 248607 236147 248641 236175
rect 248669 236147 248703 236175
rect 248731 236147 248779 236175
rect 248469 236113 248779 236147
rect 248469 236085 248517 236113
rect 248545 236085 248579 236113
rect 248607 236085 248641 236113
rect 248669 236085 248703 236113
rect 248731 236085 248779 236113
rect 248469 236051 248779 236085
rect 248469 236023 248517 236051
rect 248545 236023 248579 236051
rect 248607 236023 248641 236051
rect 248669 236023 248703 236051
rect 248731 236023 248779 236051
rect 248469 235989 248779 236023
rect 248469 235961 248517 235989
rect 248545 235961 248579 235989
rect 248607 235961 248641 235989
rect 248669 235961 248703 235989
rect 248731 235961 248779 235989
rect 248469 227175 248779 235961
rect 248469 227147 248517 227175
rect 248545 227147 248579 227175
rect 248607 227147 248641 227175
rect 248669 227147 248703 227175
rect 248731 227147 248779 227175
rect 248469 227113 248779 227147
rect 248469 227085 248517 227113
rect 248545 227085 248579 227113
rect 248607 227085 248641 227113
rect 248669 227085 248703 227113
rect 248731 227085 248779 227113
rect 248469 227051 248779 227085
rect 248469 227023 248517 227051
rect 248545 227023 248579 227051
rect 248607 227023 248641 227051
rect 248669 227023 248703 227051
rect 248731 227023 248779 227051
rect 248469 226989 248779 227023
rect 248469 226961 248517 226989
rect 248545 226961 248579 226989
rect 248607 226961 248641 226989
rect 248669 226961 248703 226989
rect 248731 226961 248779 226989
rect 248469 218175 248779 226961
rect 248469 218147 248517 218175
rect 248545 218147 248579 218175
rect 248607 218147 248641 218175
rect 248669 218147 248703 218175
rect 248731 218147 248779 218175
rect 248469 218113 248779 218147
rect 248469 218085 248517 218113
rect 248545 218085 248579 218113
rect 248607 218085 248641 218113
rect 248669 218085 248703 218113
rect 248731 218085 248779 218113
rect 248469 218051 248779 218085
rect 248469 218023 248517 218051
rect 248545 218023 248579 218051
rect 248607 218023 248641 218051
rect 248669 218023 248703 218051
rect 248731 218023 248779 218051
rect 248469 217989 248779 218023
rect 248469 217961 248517 217989
rect 248545 217961 248579 217989
rect 248607 217961 248641 217989
rect 248669 217961 248703 217989
rect 248731 217961 248779 217989
rect 248469 209175 248779 217961
rect 248469 209147 248517 209175
rect 248545 209147 248579 209175
rect 248607 209147 248641 209175
rect 248669 209147 248703 209175
rect 248731 209147 248779 209175
rect 248469 209113 248779 209147
rect 248469 209085 248517 209113
rect 248545 209085 248579 209113
rect 248607 209085 248641 209113
rect 248669 209085 248703 209113
rect 248731 209085 248779 209113
rect 248469 209051 248779 209085
rect 248469 209023 248517 209051
rect 248545 209023 248579 209051
rect 248607 209023 248641 209051
rect 248669 209023 248703 209051
rect 248731 209023 248779 209051
rect 248469 208989 248779 209023
rect 248469 208961 248517 208989
rect 248545 208961 248579 208989
rect 248607 208961 248641 208989
rect 248669 208961 248703 208989
rect 248731 208961 248779 208989
rect 248469 200175 248779 208961
rect 248469 200147 248517 200175
rect 248545 200147 248579 200175
rect 248607 200147 248641 200175
rect 248669 200147 248703 200175
rect 248731 200147 248779 200175
rect 248469 200113 248779 200147
rect 248469 200085 248517 200113
rect 248545 200085 248579 200113
rect 248607 200085 248641 200113
rect 248669 200085 248703 200113
rect 248731 200085 248779 200113
rect 248469 200051 248779 200085
rect 248469 200023 248517 200051
rect 248545 200023 248579 200051
rect 248607 200023 248641 200051
rect 248669 200023 248703 200051
rect 248731 200023 248779 200051
rect 248469 199989 248779 200023
rect 248469 199961 248517 199989
rect 248545 199961 248579 199989
rect 248607 199961 248641 199989
rect 248669 199961 248703 199989
rect 248731 199961 248779 199989
rect 248469 191175 248779 199961
rect 248469 191147 248517 191175
rect 248545 191147 248579 191175
rect 248607 191147 248641 191175
rect 248669 191147 248703 191175
rect 248731 191147 248779 191175
rect 248469 191113 248779 191147
rect 248469 191085 248517 191113
rect 248545 191085 248579 191113
rect 248607 191085 248641 191113
rect 248669 191085 248703 191113
rect 248731 191085 248779 191113
rect 248469 191051 248779 191085
rect 248469 191023 248517 191051
rect 248545 191023 248579 191051
rect 248607 191023 248641 191051
rect 248669 191023 248703 191051
rect 248731 191023 248779 191051
rect 248469 190989 248779 191023
rect 248469 190961 248517 190989
rect 248545 190961 248579 190989
rect 248607 190961 248641 190989
rect 248669 190961 248703 190989
rect 248731 190961 248779 190989
rect 248469 187679 248779 190961
rect 250329 299086 250639 299134
rect 250329 299058 250377 299086
rect 250405 299058 250439 299086
rect 250467 299058 250501 299086
rect 250529 299058 250563 299086
rect 250591 299058 250639 299086
rect 250329 299024 250639 299058
rect 250329 298996 250377 299024
rect 250405 298996 250439 299024
rect 250467 298996 250501 299024
rect 250529 298996 250563 299024
rect 250591 298996 250639 299024
rect 250329 298962 250639 298996
rect 250329 298934 250377 298962
rect 250405 298934 250439 298962
rect 250467 298934 250501 298962
rect 250529 298934 250563 298962
rect 250591 298934 250639 298962
rect 250329 298900 250639 298934
rect 250329 298872 250377 298900
rect 250405 298872 250439 298900
rect 250467 298872 250501 298900
rect 250529 298872 250563 298900
rect 250591 298872 250639 298900
rect 250329 293175 250639 298872
rect 250329 293147 250377 293175
rect 250405 293147 250439 293175
rect 250467 293147 250501 293175
rect 250529 293147 250563 293175
rect 250591 293147 250639 293175
rect 250329 293113 250639 293147
rect 250329 293085 250377 293113
rect 250405 293085 250439 293113
rect 250467 293085 250501 293113
rect 250529 293085 250563 293113
rect 250591 293085 250639 293113
rect 250329 293051 250639 293085
rect 250329 293023 250377 293051
rect 250405 293023 250439 293051
rect 250467 293023 250501 293051
rect 250529 293023 250563 293051
rect 250591 293023 250639 293051
rect 250329 292989 250639 293023
rect 250329 292961 250377 292989
rect 250405 292961 250439 292989
rect 250467 292961 250501 292989
rect 250529 292961 250563 292989
rect 250591 292961 250639 292989
rect 250329 284175 250639 292961
rect 250329 284147 250377 284175
rect 250405 284147 250439 284175
rect 250467 284147 250501 284175
rect 250529 284147 250563 284175
rect 250591 284147 250639 284175
rect 250329 284113 250639 284147
rect 250329 284085 250377 284113
rect 250405 284085 250439 284113
rect 250467 284085 250501 284113
rect 250529 284085 250563 284113
rect 250591 284085 250639 284113
rect 250329 284051 250639 284085
rect 250329 284023 250377 284051
rect 250405 284023 250439 284051
rect 250467 284023 250501 284051
rect 250529 284023 250563 284051
rect 250591 284023 250639 284051
rect 250329 283989 250639 284023
rect 250329 283961 250377 283989
rect 250405 283961 250439 283989
rect 250467 283961 250501 283989
rect 250529 283961 250563 283989
rect 250591 283961 250639 283989
rect 250329 275175 250639 283961
rect 250329 275147 250377 275175
rect 250405 275147 250439 275175
rect 250467 275147 250501 275175
rect 250529 275147 250563 275175
rect 250591 275147 250639 275175
rect 250329 275113 250639 275147
rect 250329 275085 250377 275113
rect 250405 275085 250439 275113
rect 250467 275085 250501 275113
rect 250529 275085 250563 275113
rect 250591 275085 250639 275113
rect 250329 275051 250639 275085
rect 250329 275023 250377 275051
rect 250405 275023 250439 275051
rect 250467 275023 250501 275051
rect 250529 275023 250563 275051
rect 250591 275023 250639 275051
rect 250329 274989 250639 275023
rect 250329 274961 250377 274989
rect 250405 274961 250439 274989
rect 250467 274961 250501 274989
rect 250529 274961 250563 274989
rect 250591 274961 250639 274989
rect 250329 266175 250639 274961
rect 250329 266147 250377 266175
rect 250405 266147 250439 266175
rect 250467 266147 250501 266175
rect 250529 266147 250563 266175
rect 250591 266147 250639 266175
rect 250329 266113 250639 266147
rect 250329 266085 250377 266113
rect 250405 266085 250439 266113
rect 250467 266085 250501 266113
rect 250529 266085 250563 266113
rect 250591 266085 250639 266113
rect 250329 266051 250639 266085
rect 250329 266023 250377 266051
rect 250405 266023 250439 266051
rect 250467 266023 250501 266051
rect 250529 266023 250563 266051
rect 250591 266023 250639 266051
rect 250329 265989 250639 266023
rect 250329 265961 250377 265989
rect 250405 265961 250439 265989
rect 250467 265961 250501 265989
rect 250529 265961 250563 265989
rect 250591 265961 250639 265989
rect 250329 257175 250639 265961
rect 250329 257147 250377 257175
rect 250405 257147 250439 257175
rect 250467 257147 250501 257175
rect 250529 257147 250563 257175
rect 250591 257147 250639 257175
rect 250329 257113 250639 257147
rect 250329 257085 250377 257113
rect 250405 257085 250439 257113
rect 250467 257085 250501 257113
rect 250529 257085 250563 257113
rect 250591 257085 250639 257113
rect 250329 257051 250639 257085
rect 250329 257023 250377 257051
rect 250405 257023 250439 257051
rect 250467 257023 250501 257051
rect 250529 257023 250563 257051
rect 250591 257023 250639 257051
rect 250329 256989 250639 257023
rect 250329 256961 250377 256989
rect 250405 256961 250439 256989
rect 250467 256961 250501 256989
rect 250529 256961 250563 256989
rect 250591 256961 250639 256989
rect 250329 248175 250639 256961
rect 250329 248147 250377 248175
rect 250405 248147 250439 248175
rect 250467 248147 250501 248175
rect 250529 248147 250563 248175
rect 250591 248147 250639 248175
rect 250329 248113 250639 248147
rect 250329 248085 250377 248113
rect 250405 248085 250439 248113
rect 250467 248085 250501 248113
rect 250529 248085 250563 248113
rect 250591 248085 250639 248113
rect 250329 248051 250639 248085
rect 250329 248023 250377 248051
rect 250405 248023 250439 248051
rect 250467 248023 250501 248051
rect 250529 248023 250563 248051
rect 250591 248023 250639 248051
rect 250329 247989 250639 248023
rect 250329 247961 250377 247989
rect 250405 247961 250439 247989
rect 250467 247961 250501 247989
rect 250529 247961 250563 247989
rect 250591 247961 250639 247989
rect 250329 239175 250639 247961
rect 250329 239147 250377 239175
rect 250405 239147 250439 239175
rect 250467 239147 250501 239175
rect 250529 239147 250563 239175
rect 250591 239147 250639 239175
rect 250329 239113 250639 239147
rect 250329 239085 250377 239113
rect 250405 239085 250439 239113
rect 250467 239085 250501 239113
rect 250529 239085 250563 239113
rect 250591 239085 250639 239113
rect 250329 239051 250639 239085
rect 250329 239023 250377 239051
rect 250405 239023 250439 239051
rect 250467 239023 250501 239051
rect 250529 239023 250563 239051
rect 250591 239023 250639 239051
rect 250329 238989 250639 239023
rect 250329 238961 250377 238989
rect 250405 238961 250439 238989
rect 250467 238961 250501 238989
rect 250529 238961 250563 238989
rect 250591 238961 250639 238989
rect 250329 230175 250639 238961
rect 250329 230147 250377 230175
rect 250405 230147 250439 230175
rect 250467 230147 250501 230175
rect 250529 230147 250563 230175
rect 250591 230147 250639 230175
rect 250329 230113 250639 230147
rect 250329 230085 250377 230113
rect 250405 230085 250439 230113
rect 250467 230085 250501 230113
rect 250529 230085 250563 230113
rect 250591 230085 250639 230113
rect 250329 230051 250639 230085
rect 250329 230023 250377 230051
rect 250405 230023 250439 230051
rect 250467 230023 250501 230051
rect 250529 230023 250563 230051
rect 250591 230023 250639 230051
rect 250329 229989 250639 230023
rect 250329 229961 250377 229989
rect 250405 229961 250439 229989
rect 250467 229961 250501 229989
rect 250529 229961 250563 229989
rect 250591 229961 250639 229989
rect 250329 221175 250639 229961
rect 250329 221147 250377 221175
rect 250405 221147 250439 221175
rect 250467 221147 250501 221175
rect 250529 221147 250563 221175
rect 250591 221147 250639 221175
rect 250329 221113 250639 221147
rect 250329 221085 250377 221113
rect 250405 221085 250439 221113
rect 250467 221085 250501 221113
rect 250529 221085 250563 221113
rect 250591 221085 250639 221113
rect 250329 221051 250639 221085
rect 250329 221023 250377 221051
rect 250405 221023 250439 221051
rect 250467 221023 250501 221051
rect 250529 221023 250563 221051
rect 250591 221023 250639 221051
rect 250329 220989 250639 221023
rect 250329 220961 250377 220989
rect 250405 220961 250439 220989
rect 250467 220961 250501 220989
rect 250529 220961 250563 220989
rect 250591 220961 250639 220989
rect 250329 212175 250639 220961
rect 250329 212147 250377 212175
rect 250405 212147 250439 212175
rect 250467 212147 250501 212175
rect 250529 212147 250563 212175
rect 250591 212147 250639 212175
rect 250329 212113 250639 212147
rect 250329 212085 250377 212113
rect 250405 212085 250439 212113
rect 250467 212085 250501 212113
rect 250529 212085 250563 212113
rect 250591 212085 250639 212113
rect 250329 212051 250639 212085
rect 250329 212023 250377 212051
rect 250405 212023 250439 212051
rect 250467 212023 250501 212051
rect 250529 212023 250563 212051
rect 250591 212023 250639 212051
rect 250329 211989 250639 212023
rect 250329 211961 250377 211989
rect 250405 211961 250439 211989
rect 250467 211961 250501 211989
rect 250529 211961 250563 211989
rect 250591 211961 250639 211989
rect 250329 203175 250639 211961
rect 250329 203147 250377 203175
rect 250405 203147 250439 203175
rect 250467 203147 250501 203175
rect 250529 203147 250563 203175
rect 250591 203147 250639 203175
rect 250329 203113 250639 203147
rect 250329 203085 250377 203113
rect 250405 203085 250439 203113
rect 250467 203085 250501 203113
rect 250529 203085 250563 203113
rect 250591 203085 250639 203113
rect 250329 203051 250639 203085
rect 250329 203023 250377 203051
rect 250405 203023 250439 203051
rect 250467 203023 250501 203051
rect 250529 203023 250563 203051
rect 250591 203023 250639 203051
rect 250329 202989 250639 203023
rect 250329 202961 250377 202989
rect 250405 202961 250439 202989
rect 250467 202961 250501 202989
rect 250529 202961 250563 202989
rect 250591 202961 250639 202989
rect 250329 194175 250639 202961
rect 250329 194147 250377 194175
rect 250405 194147 250439 194175
rect 250467 194147 250501 194175
rect 250529 194147 250563 194175
rect 250591 194147 250639 194175
rect 250329 194113 250639 194147
rect 250329 194085 250377 194113
rect 250405 194085 250439 194113
rect 250467 194085 250501 194113
rect 250529 194085 250563 194113
rect 250591 194085 250639 194113
rect 250329 194051 250639 194085
rect 250329 194023 250377 194051
rect 250405 194023 250439 194051
rect 250467 194023 250501 194051
rect 250529 194023 250563 194051
rect 250591 194023 250639 194051
rect 250329 193989 250639 194023
rect 250329 193961 250377 193989
rect 250405 193961 250439 193989
rect 250467 193961 250501 193989
rect 250529 193961 250563 193989
rect 250591 193961 250639 193989
rect 250329 187679 250639 193961
rect 263829 298606 264139 299134
rect 263829 298578 263877 298606
rect 263905 298578 263939 298606
rect 263967 298578 264001 298606
rect 264029 298578 264063 298606
rect 264091 298578 264139 298606
rect 263829 298544 264139 298578
rect 263829 298516 263877 298544
rect 263905 298516 263939 298544
rect 263967 298516 264001 298544
rect 264029 298516 264063 298544
rect 264091 298516 264139 298544
rect 263829 298482 264139 298516
rect 263829 298454 263877 298482
rect 263905 298454 263939 298482
rect 263967 298454 264001 298482
rect 264029 298454 264063 298482
rect 264091 298454 264139 298482
rect 263829 298420 264139 298454
rect 263829 298392 263877 298420
rect 263905 298392 263939 298420
rect 263967 298392 264001 298420
rect 264029 298392 264063 298420
rect 264091 298392 264139 298420
rect 263829 290175 264139 298392
rect 263829 290147 263877 290175
rect 263905 290147 263939 290175
rect 263967 290147 264001 290175
rect 264029 290147 264063 290175
rect 264091 290147 264139 290175
rect 263829 290113 264139 290147
rect 263829 290085 263877 290113
rect 263905 290085 263939 290113
rect 263967 290085 264001 290113
rect 264029 290085 264063 290113
rect 264091 290085 264139 290113
rect 263829 290051 264139 290085
rect 263829 290023 263877 290051
rect 263905 290023 263939 290051
rect 263967 290023 264001 290051
rect 264029 290023 264063 290051
rect 264091 290023 264139 290051
rect 263829 289989 264139 290023
rect 263829 289961 263877 289989
rect 263905 289961 263939 289989
rect 263967 289961 264001 289989
rect 264029 289961 264063 289989
rect 264091 289961 264139 289989
rect 263829 281175 264139 289961
rect 263829 281147 263877 281175
rect 263905 281147 263939 281175
rect 263967 281147 264001 281175
rect 264029 281147 264063 281175
rect 264091 281147 264139 281175
rect 263829 281113 264139 281147
rect 263829 281085 263877 281113
rect 263905 281085 263939 281113
rect 263967 281085 264001 281113
rect 264029 281085 264063 281113
rect 264091 281085 264139 281113
rect 263829 281051 264139 281085
rect 263829 281023 263877 281051
rect 263905 281023 263939 281051
rect 263967 281023 264001 281051
rect 264029 281023 264063 281051
rect 264091 281023 264139 281051
rect 263829 280989 264139 281023
rect 263829 280961 263877 280989
rect 263905 280961 263939 280989
rect 263967 280961 264001 280989
rect 264029 280961 264063 280989
rect 264091 280961 264139 280989
rect 263829 272175 264139 280961
rect 263829 272147 263877 272175
rect 263905 272147 263939 272175
rect 263967 272147 264001 272175
rect 264029 272147 264063 272175
rect 264091 272147 264139 272175
rect 263829 272113 264139 272147
rect 263829 272085 263877 272113
rect 263905 272085 263939 272113
rect 263967 272085 264001 272113
rect 264029 272085 264063 272113
rect 264091 272085 264139 272113
rect 263829 272051 264139 272085
rect 263829 272023 263877 272051
rect 263905 272023 263939 272051
rect 263967 272023 264001 272051
rect 264029 272023 264063 272051
rect 264091 272023 264139 272051
rect 263829 271989 264139 272023
rect 263829 271961 263877 271989
rect 263905 271961 263939 271989
rect 263967 271961 264001 271989
rect 264029 271961 264063 271989
rect 264091 271961 264139 271989
rect 263829 263175 264139 271961
rect 263829 263147 263877 263175
rect 263905 263147 263939 263175
rect 263967 263147 264001 263175
rect 264029 263147 264063 263175
rect 264091 263147 264139 263175
rect 263829 263113 264139 263147
rect 263829 263085 263877 263113
rect 263905 263085 263939 263113
rect 263967 263085 264001 263113
rect 264029 263085 264063 263113
rect 264091 263085 264139 263113
rect 263829 263051 264139 263085
rect 263829 263023 263877 263051
rect 263905 263023 263939 263051
rect 263967 263023 264001 263051
rect 264029 263023 264063 263051
rect 264091 263023 264139 263051
rect 263829 262989 264139 263023
rect 263829 262961 263877 262989
rect 263905 262961 263939 262989
rect 263967 262961 264001 262989
rect 264029 262961 264063 262989
rect 264091 262961 264139 262989
rect 263829 254175 264139 262961
rect 263829 254147 263877 254175
rect 263905 254147 263939 254175
rect 263967 254147 264001 254175
rect 264029 254147 264063 254175
rect 264091 254147 264139 254175
rect 263829 254113 264139 254147
rect 263829 254085 263877 254113
rect 263905 254085 263939 254113
rect 263967 254085 264001 254113
rect 264029 254085 264063 254113
rect 264091 254085 264139 254113
rect 263829 254051 264139 254085
rect 263829 254023 263877 254051
rect 263905 254023 263939 254051
rect 263967 254023 264001 254051
rect 264029 254023 264063 254051
rect 264091 254023 264139 254051
rect 263829 253989 264139 254023
rect 263829 253961 263877 253989
rect 263905 253961 263939 253989
rect 263967 253961 264001 253989
rect 264029 253961 264063 253989
rect 264091 253961 264139 253989
rect 263829 245175 264139 253961
rect 263829 245147 263877 245175
rect 263905 245147 263939 245175
rect 263967 245147 264001 245175
rect 264029 245147 264063 245175
rect 264091 245147 264139 245175
rect 263829 245113 264139 245147
rect 263829 245085 263877 245113
rect 263905 245085 263939 245113
rect 263967 245085 264001 245113
rect 264029 245085 264063 245113
rect 264091 245085 264139 245113
rect 263829 245051 264139 245085
rect 263829 245023 263877 245051
rect 263905 245023 263939 245051
rect 263967 245023 264001 245051
rect 264029 245023 264063 245051
rect 264091 245023 264139 245051
rect 263829 244989 264139 245023
rect 263829 244961 263877 244989
rect 263905 244961 263939 244989
rect 263967 244961 264001 244989
rect 264029 244961 264063 244989
rect 264091 244961 264139 244989
rect 263829 236175 264139 244961
rect 263829 236147 263877 236175
rect 263905 236147 263939 236175
rect 263967 236147 264001 236175
rect 264029 236147 264063 236175
rect 264091 236147 264139 236175
rect 263829 236113 264139 236147
rect 263829 236085 263877 236113
rect 263905 236085 263939 236113
rect 263967 236085 264001 236113
rect 264029 236085 264063 236113
rect 264091 236085 264139 236113
rect 263829 236051 264139 236085
rect 263829 236023 263877 236051
rect 263905 236023 263939 236051
rect 263967 236023 264001 236051
rect 264029 236023 264063 236051
rect 264091 236023 264139 236051
rect 263829 235989 264139 236023
rect 263829 235961 263877 235989
rect 263905 235961 263939 235989
rect 263967 235961 264001 235989
rect 264029 235961 264063 235989
rect 264091 235961 264139 235989
rect 263829 227175 264139 235961
rect 263829 227147 263877 227175
rect 263905 227147 263939 227175
rect 263967 227147 264001 227175
rect 264029 227147 264063 227175
rect 264091 227147 264139 227175
rect 263829 227113 264139 227147
rect 263829 227085 263877 227113
rect 263905 227085 263939 227113
rect 263967 227085 264001 227113
rect 264029 227085 264063 227113
rect 264091 227085 264139 227113
rect 263829 227051 264139 227085
rect 263829 227023 263877 227051
rect 263905 227023 263939 227051
rect 263967 227023 264001 227051
rect 264029 227023 264063 227051
rect 264091 227023 264139 227051
rect 263829 226989 264139 227023
rect 263829 226961 263877 226989
rect 263905 226961 263939 226989
rect 263967 226961 264001 226989
rect 264029 226961 264063 226989
rect 264091 226961 264139 226989
rect 263829 218175 264139 226961
rect 263829 218147 263877 218175
rect 263905 218147 263939 218175
rect 263967 218147 264001 218175
rect 264029 218147 264063 218175
rect 264091 218147 264139 218175
rect 263829 218113 264139 218147
rect 263829 218085 263877 218113
rect 263905 218085 263939 218113
rect 263967 218085 264001 218113
rect 264029 218085 264063 218113
rect 264091 218085 264139 218113
rect 263829 218051 264139 218085
rect 263829 218023 263877 218051
rect 263905 218023 263939 218051
rect 263967 218023 264001 218051
rect 264029 218023 264063 218051
rect 264091 218023 264139 218051
rect 263829 217989 264139 218023
rect 263829 217961 263877 217989
rect 263905 217961 263939 217989
rect 263967 217961 264001 217989
rect 264029 217961 264063 217989
rect 264091 217961 264139 217989
rect 263829 209175 264139 217961
rect 263829 209147 263877 209175
rect 263905 209147 263939 209175
rect 263967 209147 264001 209175
rect 264029 209147 264063 209175
rect 264091 209147 264139 209175
rect 263829 209113 264139 209147
rect 263829 209085 263877 209113
rect 263905 209085 263939 209113
rect 263967 209085 264001 209113
rect 264029 209085 264063 209113
rect 264091 209085 264139 209113
rect 263829 209051 264139 209085
rect 263829 209023 263877 209051
rect 263905 209023 263939 209051
rect 263967 209023 264001 209051
rect 264029 209023 264063 209051
rect 264091 209023 264139 209051
rect 263829 208989 264139 209023
rect 263829 208961 263877 208989
rect 263905 208961 263939 208989
rect 263967 208961 264001 208989
rect 264029 208961 264063 208989
rect 264091 208961 264139 208989
rect 263829 200175 264139 208961
rect 263829 200147 263877 200175
rect 263905 200147 263939 200175
rect 263967 200147 264001 200175
rect 264029 200147 264063 200175
rect 264091 200147 264139 200175
rect 263829 200113 264139 200147
rect 263829 200085 263877 200113
rect 263905 200085 263939 200113
rect 263967 200085 264001 200113
rect 264029 200085 264063 200113
rect 264091 200085 264139 200113
rect 263829 200051 264139 200085
rect 263829 200023 263877 200051
rect 263905 200023 263939 200051
rect 263967 200023 264001 200051
rect 264029 200023 264063 200051
rect 264091 200023 264139 200051
rect 263829 199989 264139 200023
rect 263829 199961 263877 199989
rect 263905 199961 263939 199989
rect 263967 199961 264001 199989
rect 264029 199961 264063 199989
rect 264091 199961 264139 199989
rect 263829 191175 264139 199961
rect 263829 191147 263877 191175
rect 263905 191147 263939 191175
rect 263967 191147 264001 191175
rect 264029 191147 264063 191175
rect 264091 191147 264139 191175
rect 263829 191113 264139 191147
rect 263829 191085 263877 191113
rect 263905 191085 263939 191113
rect 263967 191085 264001 191113
rect 264029 191085 264063 191113
rect 264091 191085 264139 191113
rect 263829 191051 264139 191085
rect 263829 191023 263877 191051
rect 263905 191023 263939 191051
rect 263967 191023 264001 191051
rect 264029 191023 264063 191051
rect 264091 191023 264139 191051
rect 263829 190989 264139 191023
rect 263829 190961 263877 190989
rect 263905 190961 263939 190989
rect 263967 190961 264001 190989
rect 264029 190961 264063 190989
rect 264091 190961 264139 190989
rect 234969 185147 235017 185175
rect 235045 185147 235079 185175
rect 235107 185147 235141 185175
rect 235169 185147 235203 185175
rect 235231 185147 235279 185175
rect 234969 185113 235279 185147
rect 234969 185085 235017 185113
rect 235045 185085 235079 185113
rect 235107 185085 235141 185113
rect 235169 185085 235203 185113
rect 235231 185085 235279 185113
rect 234969 185051 235279 185085
rect 234969 185023 235017 185051
rect 235045 185023 235079 185051
rect 235107 185023 235141 185051
rect 235169 185023 235203 185051
rect 235231 185023 235279 185051
rect 234969 184989 235279 185023
rect 234969 184961 235017 184989
rect 235045 184961 235079 184989
rect 235107 184961 235141 184989
rect 235169 184961 235203 184989
rect 235231 184961 235279 184989
rect 234969 176175 235279 184961
rect 244904 185175 245064 185192
rect 244904 185147 244939 185175
rect 244967 185147 245001 185175
rect 245029 185147 245064 185175
rect 244904 185113 245064 185147
rect 244904 185085 244939 185113
rect 244967 185085 245001 185113
rect 245029 185085 245064 185113
rect 244904 185051 245064 185085
rect 244904 185023 244939 185051
rect 244967 185023 245001 185051
rect 245029 185023 245064 185051
rect 244904 184989 245064 185023
rect 244904 184961 244939 184989
rect 244967 184961 245001 184989
rect 245029 184961 245064 184989
rect 244904 184944 245064 184961
rect 237224 182175 237384 182192
rect 237224 182147 237259 182175
rect 237287 182147 237321 182175
rect 237349 182147 237384 182175
rect 237224 182113 237384 182147
rect 237224 182085 237259 182113
rect 237287 182085 237321 182113
rect 237349 182085 237384 182113
rect 237224 182051 237384 182085
rect 237224 182023 237259 182051
rect 237287 182023 237321 182051
rect 237349 182023 237384 182051
rect 237224 181989 237384 182023
rect 237224 181961 237259 181989
rect 237287 181961 237321 181989
rect 237349 181961 237384 181989
rect 237224 181944 237384 181961
rect 252584 182175 252744 182192
rect 252584 182147 252619 182175
rect 252647 182147 252681 182175
rect 252709 182147 252744 182175
rect 252584 182113 252744 182147
rect 252584 182085 252619 182113
rect 252647 182085 252681 182113
rect 252709 182085 252744 182113
rect 252584 182051 252744 182085
rect 252584 182023 252619 182051
rect 252647 182023 252681 182051
rect 252709 182023 252744 182051
rect 252584 181989 252744 182023
rect 252584 181961 252619 181989
rect 252647 181961 252681 181989
rect 252709 181961 252744 181989
rect 252584 181944 252744 181961
rect 263829 182175 264139 190961
rect 263829 182147 263877 182175
rect 263905 182147 263939 182175
rect 263967 182147 264001 182175
rect 264029 182147 264063 182175
rect 264091 182147 264139 182175
rect 263829 182113 264139 182147
rect 263829 182085 263877 182113
rect 263905 182085 263939 182113
rect 263967 182085 264001 182113
rect 264029 182085 264063 182113
rect 264091 182085 264139 182113
rect 263829 182051 264139 182085
rect 263829 182023 263877 182051
rect 263905 182023 263939 182051
rect 263967 182023 264001 182051
rect 264029 182023 264063 182051
rect 264091 182023 264139 182051
rect 263829 181989 264139 182023
rect 263829 181961 263877 181989
rect 263905 181961 263939 181989
rect 263967 181961 264001 181989
rect 264029 181961 264063 181989
rect 264091 181961 264139 181989
rect 234969 176147 235017 176175
rect 235045 176147 235079 176175
rect 235107 176147 235141 176175
rect 235169 176147 235203 176175
rect 235231 176147 235279 176175
rect 234969 176113 235279 176147
rect 234969 176085 235017 176113
rect 235045 176085 235079 176113
rect 235107 176085 235141 176113
rect 235169 176085 235203 176113
rect 235231 176085 235279 176113
rect 234969 176051 235279 176085
rect 234969 176023 235017 176051
rect 235045 176023 235079 176051
rect 235107 176023 235141 176051
rect 235169 176023 235203 176051
rect 235231 176023 235279 176051
rect 234969 175989 235279 176023
rect 234969 175961 235017 175989
rect 235045 175961 235079 175989
rect 235107 175961 235141 175989
rect 235169 175961 235203 175989
rect 235231 175961 235279 175989
rect 234969 167175 235279 175961
rect 244904 176175 245064 176192
rect 244904 176147 244939 176175
rect 244967 176147 245001 176175
rect 245029 176147 245064 176175
rect 244904 176113 245064 176147
rect 244904 176085 244939 176113
rect 244967 176085 245001 176113
rect 245029 176085 245064 176113
rect 244904 176051 245064 176085
rect 244904 176023 244939 176051
rect 244967 176023 245001 176051
rect 245029 176023 245064 176051
rect 244904 175989 245064 176023
rect 244904 175961 244939 175989
rect 244967 175961 245001 175989
rect 245029 175961 245064 175989
rect 244904 175944 245064 175961
rect 237224 173175 237384 173192
rect 237224 173147 237259 173175
rect 237287 173147 237321 173175
rect 237349 173147 237384 173175
rect 237224 173113 237384 173147
rect 237224 173085 237259 173113
rect 237287 173085 237321 173113
rect 237349 173085 237384 173113
rect 237224 173051 237384 173085
rect 237224 173023 237259 173051
rect 237287 173023 237321 173051
rect 237349 173023 237384 173051
rect 237224 172989 237384 173023
rect 237224 172961 237259 172989
rect 237287 172961 237321 172989
rect 237349 172961 237384 172989
rect 237224 172944 237384 172961
rect 252584 173175 252744 173192
rect 252584 173147 252619 173175
rect 252647 173147 252681 173175
rect 252709 173147 252744 173175
rect 252584 173113 252744 173147
rect 252584 173085 252619 173113
rect 252647 173085 252681 173113
rect 252709 173085 252744 173113
rect 252584 173051 252744 173085
rect 252584 173023 252619 173051
rect 252647 173023 252681 173051
rect 252709 173023 252744 173051
rect 252584 172989 252744 173023
rect 252584 172961 252619 172989
rect 252647 172961 252681 172989
rect 252709 172961 252744 172989
rect 252584 172944 252744 172961
rect 263829 173175 264139 181961
rect 263829 173147 263877 173175
rect 263905 173147 263939 173175
rect 263967 173147 264001 173175
rect 264029 173147 264063 173175
rect 264091 173147 264139 173175
rect 263829 173113 264139 173147
rect 263829 173085 263877 173113
rect 263905 173085 263939 173113
rect 263967 173085 264001 173113
rect 264029 173085 264063 173113
rect 264091 173085 264139 173113
rect 263829 173051 264139 173085
rect 263829 173023 263877 173051
rect 263905 173023 263939 173051
rect 263967 173023 264001 173051
rect 264029 173023 264063 173051
rect 264091 173023 264139 173051
rect 263829 172989 264139 173023
rect 263829 172961 263877 172989
rect 263905 172961 263939 172989
rect 263967 172961 264001 172989
rect 264029 172961 264063 172989
rect 264091 172961 264139 172989
rect 234969 167147 235017 167175
rect 235045 167147 235079 167175
rect 235107 167147 235141 167175
rect 235169 167147 235203 167175
rect 235231 167147 235279 167175
rect 234969 167113 235279 167147
rect 234969 167085 235017 167113
rect 235045 167085 235079 167113
rect 235107 167085 235141 167113
rect 235169 167085 235203 167113
rect 235231 167085 235279 167113
rect 234969 167051 235279 167085
rect 234969 167023 235017 167051
rect 235045 167023 235079 167051
rect 235107 167023 235141 167051
rect 235169 167023 235203 167051
rect 235231 167023 235279 167051
rect 234969 166989 235279 167023
rect 234969 166961 235017 166989
rect 235045 166961 235079 166989
rect 235107 166961 235141 166989
rect 235169 166961 235203 166989
rect 235231 166961 235279 166989
rect 234969 158175 235279 166961
rect 248469 164175 248779 172089
rect 248469 164147 248517 164175
rect 248545 164147 248579 164175
rect 248607 164147 248641 164175
rect 248669 164147 248703 164175
rect 248731 164147 248779 164175
rect 248469 164113 248779 164147
rect 248469 164085 248517 164113
rect 248545 164085 248579 164113
rect 248607 164085 248641 164113
rect 248669 164085 248703 164113
rect 248731 164085 248779 164113
rect 248469 164051 248779 164085
rect 248469 164023 248517 164051
rect 248545 164023 248579 164051
rect 248607 164023 248641 164051
rect 248669 164023 248703 164051
rect 248731 164023 248779 164051
rect 248469 163989 248779 164023
rect 248469 163961 248517 163989
rect 248545 163961 248579 163989
rect 248607 163961 248641 163989
rect 248669 163961 248703 163989
rect 248731 163961 248779 163989
rect 234969 158147 235017 158175
rect 235045 158147 235079 158175
rect 235107 158147 235141 158175
rect 235169 158147 235203 158175
rect 235231 158147 235279 158175
rect 234969 158113 235279 158147
rect 234969 158085 235017 158113
rect 235045 158085 235079 158113
rect 235107 158085 235141 158113
rect 235169 158085 235203 158113
rect 235231 158085 235279 158113
rect 234969 158051 235279 158085
rect 234969 158023 235017 158051
rect 235045 158023 235079 158051
rect 235107 158023 235141 158051
rect 235169 158023 235203 158051
rect 235231 158023 235279 158051
rect 234969 157989 235279 158023
rect 234969 157961 235017 157989
rect 235045 157961 235079 157989
rect 235107 157961 235141 157989
rect 235169 157961 235203 157989
rect 235231 157961 235279 157989
rect 234969 149175 235279 157961
rect 239584 158175 239744 158192
rect 239584 158147 239619 158175
rect 239647 158147 239681 158175
rect 239709 158147 239744 158175
rect 239584 158113 239744 158147
rect 239584 158085 239619 158113
rect 239647 158085 239681 158113
rect 239709 158085 239744 158113
rect 239584 158051 239744 158085
rect 239584 158023 239619 158051
rect 239647 158023 239681 158051
rect 239709 158023 239744 158051
rect 239584 157989 239744 158023
rect 239584 157961 239619 157989
rect 239647 157961 239681 157989
rect 239709 157961 239744 157989
rect 239584 157944 239744 157961
rect 247264 155175 247424 155192
rect 247264 155147 247299 155175
rect 247327 155147 247361 155175
rect 247389 155147 247424 155175
rect 247264 155113 247424 155147
rect 247264 155085 247299 155113
rect 247327 155085 247361 155113
rect 247389 155085 247424 155113
rect 247264 155051 247424 155085
rect 247264 155023 247299 155051
rect 247327 155023 247361 155051
rect 247389 155023 247424 155051
rect 247264 154989 247424 155023
rect 247264 154961 247299 154989
rect 247327 154961 247361 154989
rect 247389 154961 247424 154989
rect 247264 154944 247424 154961
rect 248469 155175 248779 163961
rect 248469 155147 248517 155175
rect 248545 155147 248579 155175
rect 248607 155147 248641 155175
rect 248669 155147 248703 155175
rect 248731 155147 248779 155175
rect 248469 155113 248779 155147
rect 248469 155085 248517 155113
rect 248545 155085 248579 155113
rect 248607 155085 248641 155113
rect 248669 155085 248703 155113
rect 248731 155085 248779 155113
rect 248469 155051 248779 155085
rect 248469 155023 248517 155051
rect 248545 155023 248579 155051
rect 248607 155023 248641 155051
rect 248669 155023 248703 155051
rect 248731 155023 248779 155051
rect 248469 154989 248779 155023
rect 248469 154961 248517 154989
rect 248545 154961 248579 154989
rect 248607 154961 248641 154989
rect 248669 154961 248703 154989
rect 248731 154961 248779 154989
rect 234969 149147 235017 149175
rect 235045 149147 235079 149175
rect 235107 149147 235141 149175
rect 235169 149147 235203 149175
rect 235231 149147 235279 149175
rect 234969 149113 235279 149147
rect 234969 149085 235017 149113
rect 235045 149085 235079 149113
rect 235107 149085 235141 149113
rect 235169 149085 235203 149113
rect 235231 149085 235279 149113
rect 234969 149051 235279 149085
rect 234969 149023 235017 149051
rect 235045 149023 235079 149051
rect 235107 149023 235141 149051
rect 235169 149023 235203 149051
rect 235231 149023 235279 149051
rect 234969 148989 235279 149023
rect 234969 148961 235017 148989
rect 235045 148961 235079 148989
rect 235107 148961 235141 148989
rect 235169 148961 235203 148989
rect 235231 148961 235279 148989
rect 234969 140175 235279 148961
rect 239584 149175 239744 149192
rect 239584 149147 239619 149175
rect 239647 149147 239681 149175
rect 239709 149147 239744 149175
rect 239584 149113 239744 149147
rect 239584 149085 239619 149113
rect 239647 149085 239681 149113
rect 239709 149085 239744 149113
rect 239584 149051 239744 149085
rect 239584 149023 239619 149051
rect 239647 149023 239681 149051
rect 239709 149023 239744 149051
rect 239584 148989 239744 149023
rect 239584 148961 239619 148989
rect 239647 148961 239681 148989
rect 239709 148961 239744 148989
rect 239584 148944 239744 148961
rect 247264 146175 247424 146192
rect 247264 146147 247299 146175
rect 247327 146147 247361 146175
rect 247389 146147 247424 146175
rect 247264 146113 247424 146147
rect 247264 146085 247299 146113
rect 247327 146085 247361 146113
rect 247389 146085 247424 146113
rect 247264 146051 247424 146085
rect 247264 146023 247299 146051
rect 247327 146023 247361 146051
rect 247389 146023 247424 146051
rect 247264 145989 247424 146023
rect 247264 145961 247299 145989
rect 247327 145961 247361 145989
rect 247389 145961 247424 145989
rect 247264 145944 247424 145961
rect 248469 146175 248779 154961
rect 248469 146147 248517 146175
rect 248545 146147 248579 146175
rect 248607 146147 248641 146175
rect 248669 146147 248703 146175
rect 248731 146147 248779 146175
rect 248469 146113 248779 146147
rect 248469 146085 248517 146113
rect 248545 146085 248579 146113
rect 248607 146085 248641 146113
rect 248669 146085 248703 146113
rect 248731 146085 248779 146113
rect 248469 146051 248779 146085
rect 248469 146023 248517 146051
rect 248545 146023 248579 146051
rect 248607 146023 248641 146051
rect 248669 146023 248703 146051
rect 248731 146023 248779 146051
rect 248469 145989 248779 146023
rect 248469 145961 248517 145989
rect 248545 145961 248579 145989
rect 248607 145961 248641 145989
rect 248669 145961 248703 145989
rect 248731 145961 248779 145989
rect 234969 140147 235017 140175
rect 235045 140147 235079 140175
rect 235107 140147 235141 140175
rect 235169 140147 235203 140175
rect 235231 140147 235279 140175
rect 234969 140113 235279 140147
rect 234969 140085 235017 140113
rect 235045 140085 235079 140113
rect 235107 140085 235141 140113
rect 235169 140085 235203 140113
rect 235231 140085 235279 140113
rect 234969 140051 235279 140085
rect 234969 140023 235017 140051
rect 235045 140023 235079 140051
rect 235107 140023 235141 140051
rect 235169 140023 235203 140051
rect 235231 140023 235279 140051
rect 234969 139989 235279 140023
rect 234969 139961 235017 139989
rect 235045 139961 235079 139989
rect 235107 139961 235141 139989
rect 235169 139961 235203 139989
rect 235231 139961 235279 139989
rect 234969 131175 235279 139961
rect 239584 140175 239744 140192
rect 239584 140147 239619 140175
rect 239647 140147 239681 140175
rect 239709 140147 239744 140175
rect 239584 140113 239744 140147
rect 239584 140085 239619 140113
rect 239647 140085 239681 140113
rect 239709 140085 239744 140113
rect 239584 140051 239744 140085
rect 239584 140023 239619 140051
rect 239647 140023 239681 140051
rect 239709 140023 239744 140051
rect 239584 139989 239744 140023
rect 239584 139961 239619 139989
rect 239647 139961 239681 139989
rect 239709 139961 239744 139989
rect 239584 139944 239744 139961
rect 247264 137175 247424 137192
rect 247264 137147 247299 137175
rect 247327 137147 247361 137175
rect 247389 137147 247424 137175
rect 247264 137113 247424 137147
rect 247264 137085 247299 137113
rect 247327 137085 247361 137113
rect 247389 137085 247424 137113
rect 247264 137051 247424 137085
rect 247264 137023 247299 137051
rect 247327 137023 247361 137051
rect 247389 137023 247424 137051
rect 247264 136989 247424 137023
rect 247264 136961 247299 136989
rect 247327 136961 247361 136989
rect 247389 136961 247424 136989
rect 247264 136944 247424 136961
rect 248469 137175 248779 145961
rect 248469 137147 248517 137175
rect 248545 137147 248579 137175
rect 248607 137147 248641 137175
rect 248669 137147 248703 137175
rect 248731 137147 248779 137175
rect 248469 137113 248779 137147
rect 248469 137085 248517 137113
rect 248545 137085 248579 137113
rect 248607 137085 248641 137113
rect 248669 137085 248703 137113
rect 248731 137085 248779 137113
rect 248469 137051 248779 137085
rect 248469 137023 248517 137051
rect 248545 137023 248579 137051
rect 248607 137023 248641 137051
rect 248669 137023 248703 137051
rect 248731 137023 248779 137051
rect 248469 136989 248779 137023
rect 248469 136961 248517 136989
rect 248545 136961 248579 136989
rect 248607 136961 248641 136989
rect 248669 136961 248703 136989
rect 248731 136961 248779 136989
rect 234969 131147 235017 131175
rect 235045 131147 235079 131175
rect 235107 131147 235141 131175
rect 235169 131147 235203 131175
rect 235231 131147 235279 131175
rect 234969 131113 235279 131147
rect 234969 131085 235017 131113
rect 235045 131085 235079 131113
rect 235107 131085 235141 131113
rect 235169 131085 235203 131113
rect 235231 131085 235279 131113
rect 234969 131051 235279 131085
rect 234969 131023 235017 131051
rect 235045 131023 235079 131051
rect 235107 131023 235141 131051
rect 235169 131023 235203 131051
rect 235231 131023 235279 131051
rect 234969 130989 235279 131023
rect 234969 130961 235017 130989
rect 235045 130961 235079 130989
rect 235107 130961 235141 130989
rect 235169 130961 235203 130989
rect 235231 130961 235279 130989
rect 234969 125367 235279 130961
rect 248469 128175 248779 136961
rect 248469 128147 248517 128175
rect 248545 128147 248579 128175
rect 248607 128147 248641 128175
rect 248669 128147 248703 128175
rect 248731 128147 248779 128175
rect 248469 128113 248779 128147
rect 248469 128085 248517 128113
rect 248545 128085 248579 128113
rect 248607 128085 248641 128113
rect 248669 128085 248703 128113
rect 248731 128085 248779 128113
rect 248469 128051 248779 128085
rect 248469 128023 248517 128051
rect 248545 128023 248579 128051
rect 248607 128023 248641 128051
rect 248669 128023 248703 128051
rect 248731 128023 248779 128051
rect 248469 127989 248779 128023
rect 248469 127961 248517 127989
rect 248545 127961 248579 127989
rect 248607 127961 248641 127989
rect 248669 127961 248703 127989
rect 248731 127961 248779 127989
rect 248469 125367 248779 127961
rect 250329 167175 250639 172089
rect 250329 167147 250377 167175
rect 250405 167147 250439 167175
rect 250467 167147 250501 167175
rect 250529 167147 250563 167175
rect 250591 167147 250639 167175
rect 250329 167113 250639 167147
rect 250329 167085 250377 167113
rect 250405 167085 250439 167113
rect 250467 167085 250501 167113
rect 250529 167085 250563 167113
rect 250591 167085 250639 167113
rect 250329 167051 250639 167085
rect 250329 167023 250377 167051
rect 250405 167023 250439 167051
rect 250467 167023 250501 167051
rect 250529 167023 250563 167051
rect 250591 167023 250639 167051
rect 250329 166989 250639 167023
rect 250329 166961 250377 166989
rect 250405 166961 250439 166989
rect 250467 166961 250501 166989
rect 250529 166961 250563 166989
rect 250591 166961 250639 166989
rect 250329 158175 250639 166961
rect 263829 164175 264139 172961
rect 263829 164147 263877 164175
rect 263905 164147 263939 164175
rect 263967 164147 264001 164175
rect 264029 164147 264063 164175
rect 264091 164147 264139 164175
rect 263829 164113 264139 164147
rect 263829 164085 263877 164113
rect 263905 164085 263939 164113
rect 263967 164085 264001 164113
rect 264029 164085 264063 164113
rect 264091 164085 264139 164113
rect 263829 164051 264139 164085
rect 263829 164023 263877 164051
rect 263905 164023 263939 164051
rect 263967 164023 264001 164051
rect 264029 164023 264063 164051
rect 264091 164023 264139 164051
rect 263829 163989 264139 164023
rect 263829 163961 263877 163989
rect 263905 163961 263939 163989
rect 263967 163961 264001 163989
rect 264029 163961 264063 163989
rect 264091 163961 264139 163989
rect 250329 158147 250377 158175
rect 250405 158147 250439 158175
rect 250467 158147 250501 158175
rect 250529 158147 250563 158175
rect 250591 158147 250639 158175
rect 250329 158113 250639 158147
rect 250329 158085 250377 158113
rect 250405 158085 250439 158113
rect 250467 158085 250501 158113
rect 250529 158085 250563 158113
rect 250591 158085 250639 158113
rect 250329 158051 250639 158085
rect 250329 158023 250377 158051
rect 250405 158023 250439 158051
rect 250467 158023 250501 158051
rect 250529 158023 250563 158051
rect 250591 158023 250639 158051
rect 250329 157989 250639 158023
rect 250329 157961 250377 157989
rect 250405 157961 250439 157989
rect 250467 157961 250501 157989
rect 250529 157961 250563 157989
rect 250591 157961 250639 157989
rect 250329 149175 250639 157961
rect 254944 158175 255104 158192
rect 254944 158147 254979 158175
rect 255007 158147 255041 158175
rect 255069 158147 255104 158175
rect 254944 158113 255104 158147
rect 254944 158085 254979 158113
rect 255007 158085 255041 158113
rect 255069 158085 255104 158113
rect 254944 158051 255104 158085
rect 254944 158023 254979 158051
rect 255007 158023 255041 158051
rect 255069 158023 255104 158051
rect 254944 157989 255104 158023
rect 254944 157961 254979 157989
rect 255007 157961 255041 157989
rect 255069 157961 255104 157989
rect 254944 157944 255104 157961
rect 262624 155175 262784 155192
rect 262624 155147 262659 155175
rect 262687 155147 262721 155175
rect 262749 155147 262784 155175
rect 262624 155113 262784 155147
rect 262624 155085 262659 155113
rect 262687 155085 262721 155113
rect 262749 155085 262784 155113
rect 262624 155051 262784 155085
rect 262624 155023 262659 155051
rect 262687 155023 262721 155051
rect 262749 155023 262784 155051
rect 262624 154989 262784 155023
rect 262624 154961 262659 154989
rect 262687 154961 262721 154989
rect 262749 154961 262784 154989
rect 262624 154944 262784 154961
rect 263829 155175 264139 163961
rect 263829 155147 263877 155175
rect 263905 155147 263939 155175
rect 263967 155147 264001 155175
rect 264029 155147 264063 155175
rect 264091 155147 264139 155175
rect 263829 155113 264139 155147
rect 263829 155085 263877 155113
rect 263905 155085 263939 155113
rect 263967 155085 264001 155113
rect 264029 155085 264063 155113
rect 264091 155085 264139 155113
rect 263829 155051 264139 155085
rect 263829 155023 263877 155051
rect 263905 155023 263939 155051
rect 263967 155023 264001 155051
rect 264029 155023 264063 155051
rect 264091 155023 264139 155051
rect 263829 154989 264139 155023
rect 263829 154961 263877 154989
rect 263905 154961 263939 154989
rect 263967 154961 264001 154989
rect 264029 154961 264063 154989
rect 264091 154961 264139 154989
rect 250329 149147 250377 149175
rect 250405 149147 250439 149175
rect 250467 149147 250501 149175
rect 250529 149147 250563 149175
rect 250591 149147 250639 149175
rect 250329 149113 250639 149147
rect 250329 149085 250377 149113
rect 250405 149085 250439 149113
rect 250467 149085 250501 149113
rect 250529 149085 250563 149113
rect 250591 149085 250639 149113
rect 250329 149051 250639 149085
rect 250329 149023 250377 149051
rect 250405 149023 250439 149051
rect 250467 149023 250501 149051
rect 250529 149023 250563 149051
rect 250591 149023 250639 149051
rect 250329 148989 250639 149023
rect 250329 148961 250377 148989
rect 250405 148961 250439 148989
rect 250467 148961 250501 148989
rect 250529 148961 250563 148989
rect 250591 148961 250639 148989
rect 250329 140175 250639 148961
rect 254944 149175 255104 149192
rect 254944 149147 254979 149175
rect 255007 149147 255041 149175
rect 255069 149147 255104 149175
rect 254944 149113 255104 149147
rect 254944 149085 254979 149113
rect 255007 149085 255041 149113
rect 255069 149085 255104 149113
rect 254944 149051 255104 149085
rect 254944 149023 254979 149051
rect 255007 149023 255041 149051
rect 255069 149023 255104 149051
rect 254944 148989 255104 149023
rect 254944 148961 254979 148989
rect 255007 148961 255041 148989
rect 255069 148961 255104 148989
rect 254944 148944 255104 148961
rect 262624 146175 262784 146192
rect 262624 146147 262659 146175
rect 262687 146147 262721 146175
rect 262749 146147 262784 146175
rect 262624 146113 262784 146147
rect 262624 146085 262659 146113
rect 262687 146085 262721 146113
rect 262749 146085 262784 146113
rect 262624 146051 262784 146085
rect 262624 146023 262659 146051
rect 262687 146023 262721 146051
rect 262749 146023 262784 146051
rect 262624 145989 262784 146023
rect 262624 145961 262659 145989
rect 262687 145961 262721 145989
rect 262749 145961 262784 145989
rect 262624 145944 262784 145961
rect 263829 146175 264139 154961
rect 263829 146147 263877 146175
rect 263905 146147 263939 146175
rect 263967 146147 264001 146175
rect 264029 146147 264063 146175
rect 264091 146147 264139 146175
rect 263829 146113 264139 146147
rect 263829 146085 263877 146113
rect 263905 146085 263939 146113
rect 263967 146085 264001 146113
rect 264029 146085 264063 146113
rect 264091 146085 264139 146113
rect 263829 146051 264139 146085
rect 263829 146023 263877 146051
rect 263905 146023 263939 146051
rect 263967 146023 264001 146051
rect 264029 146023 264063 146051
rect 264091 146023 264139 146051
rect 263829 145989 264139 146023
rect 263829 145961 263877 145989
rect 263905 145961 263939 145989
rect 263967 145961 264001 145989
rect 264029 145961 264063 145989
rect 264091 145961 264139 145989
rect 250329 140147 250377 140175
rect 250405 140147 250439 140175
rect 250467 140147 250501 140175
rect 250529 140147 250563 140175
rect 250591 140147 250639 140175
rect 250329 140113 250639 140147
rect 250329 140085 250377 140113
rect 250405 140085 250439 140113
rect 250467 140085 250501 140113
rect 250529 140085 250563 140113
rect 250591 140085 250639 140113
rect 250329 140051 250639 140085
rect 250329 140023 250377 140051
rect 250405 140023 250439 140051
rect 250467 140023 250501 140051
rect 250529 140023 250563 140051
rect 250591 140023 250639 140051
rect 250329 139989 250639 140023
rect 250329 139961 250377 139989
rect 250405 139961 250439 139989
rect 250467 139961 250501 139989
rect 250529 139961 250563 139989
rect 250591 139961 250639 139989
rect 250329 131175 250639 139961
rect 254944 140175 255104 140192
rect 254944 140147 254979 140175
rect 255007 140147 255041 140175
rect 255069 140147 255104 140175
rect 254944 140113 255104 140147
rect 254944 140085 254979 140113
rect 255007 140085 255041 140113
rect 255069 140085 255104 140113
rect 254944 140051 255104 140085
rect 254944 140023 254979 140051
rect 255007 140023 255041 140051
rect 255069 140023 255104 140051
rect 254944 139989 255104 140023
rect 254944 139961 254979 139989
rect 255007 139961 255041 139989
rect 255069 139961 255104 139989
rect 254944 139944 255104 139961
rect 262624 137175 262784 137192
rect 262624 137147 262659 137175
rect 262687 137147 262721 137175
rect 262749 137147 262784 137175
rect 262624 137113 262784 137147
rect 262624 137085 262659 137113
rect 262687 137085 262721 137113
rect 262749 137085 262784 137113
rect 262624 137051 262784 137085
rect 262624 137023 262659 137051
rect 262687 137023 262721 137051
rect 262749 137023 262784 137051
rect 262624 136989 262784 137023
rect 262624 136961 262659 136989
rect 262687 136961 262721 136989
rect 262749 136961 262784 136989
rect 262624 136944 262784 136961
rect 263829 137175 264139 145961
rect 263829 137147 263877 137175
rect 263905 137147 263939 137175
rect 263967 137147 264001 137175
rect 264029 137147 264063 137175
rect 264091 137147 264139 137175
rect 263829 137113 264139 137147
rect 263829 137085 263877 137113
rect 263905 137085 263939 137113
rect 263967 137085 264001 137113
rect 264029 137085 264063 137113
rect 264091 137085 264139 137113
rect 263829 137051 264139 137085
rect 263829 137023 263877 137051
rect 263905 137023 263939 137051
rect 263967 137023 264001 137051
rect 264029 137023 264063 137051
rect 264091 137023 264139 137051
rect 263829 136989 264139 137023
rect 263829 136961 263877 136989
rect 263905 136961 263939 136989
rect 263967 136961 264001 136989
rect 264029 136961 264063 136989
rect 264091 136961 264139 136989
rect 250329 131147 250377 131175
rect 250405 131147 250439 131175
rect 250467 131147 250501 131175
rect 250529 131147 250563 131175
rect 250591 131147 250639 131175
rect 250329 131113 250639 131147
rect 250329 131085 250377 131113
rect 250405 131085 250439 131113
rect 250467 131085 250501 131113
rect 250529 131085 250563 131113
rect 250591 131085 250639 131113
rect 250329 131051 250639 131085
rect 250329 131023 250377 131051
rect 250405 131023 250439 131051
rect 250467 131023 250501 131051
rect 250529 131023 250563 131051
rect 250591 131023 250639 131051
rect 250329 130989 250639 131023
rect 250329 130961 250377 130989
rect 250405 130961 250439 130989
rect 250467 130961 250501 130989
rect 250529 130961 250563 130989
rect 250591 130961 250639 130989
rect 250329 125367 250639 130961
rect 263829 128175 264139 136961
rect 263829 128147 263877 128175
rect 263905 128147 263939 128175
rect 263967 128147 264001 128175
rect 264029 128147 264063 128175
rect 264091 128147 264139 128175
rect 263829 128113 264139 128147
rect 263829 128085 263877 128113
rect 263905 128085 263939 128113
rect 263967 128085 264001 128113
rect 264029 128085 264063 128113
rect 264091 128085 264139 128113
rect 263829 128051 264139 128085
rect 263829 128023 263877 128051
rect 263905 128023 263939 128051
rect 263967 128023 264001 128051
rect 264029 128023 264063 128051
rect 264091 128023 264139 128051
rect 263829 127989 264139 128023
rect 263829 127961 263877 127989
rect 263905 127961 263939 127989
rect 263967 127961 264001 127989
rect 264029 127961 264063 127989
rect 264091 127961 264139 127989
rect 263829 125367 264139 127961
rect 265689 299086 265999 299134
rect 265689 299058 265737 299086
rect 265765 299058 265799 299086
rect 265827 299058 265861 299086
rect 265889 299058 265923 299086
rect 265951 299058 265999 299086
rect 265689 299024 265999 299058
rect 265689 298996 265737 299024
rect 265765 298996 265799 299024
rect 265827 298996 265861 299024
rect 265889 298996 265923 299024
rect 265951 298996 265999 299024
rect 265689 298962 265999 298996
rect 265689 298934 265737 298962
rect 265765 298934 265799 298962
rect 265827 298934 265861 298962
rect 265889 298934 265923 298962
rect 265951 298934 265999 298962
rect 265689 298900 265999 298934
rect 265689 298872 265737 298900
rect 265765 298872 265799 298900
rect 265827 298872 265861 298900
rect 265889 298872 265923 298900
rect 265951 298872 265999 298900
rect 265689 293175 265999 298872
rect 279189 298606 279499 299134
rect 279189 298578 279237 298606
rect 279265 298578 279299 298606
rect 279327 298578 279361 298606
rect 279389 298578 279423 298606
rect 279451 298578 279499 298606
rect 279189 298544 279499 298578
rect 279189 298516 279237 298544
rect 279265 298516 279299 298544
rect 279327 298516 279361 298544
rect 279389 298516 279423 298544
rect 279451 298516 279499 298544
rect 279189 298482 279499 298516
rect 279189 298454 279237 298482
rect 279265 298454 279299 298482
rect 279327 298454 279361 298482
rect 279389 298454 279423 298482
rect 279451 298454 279499 298482
rect 279189 298420 279499 298454
rect 279189 298392 279237 298420
rect 279265 298392 279299 298420
rect 279327 298392 279361 298420
rect 279389 298392 279423 298420
rect 279451 298392 279499 298420
rect 265689 293147 265737 293175
rect 265765 293147 265799 293175
rect 265827 293147 265861 293175
rect 265889 293147 265923 293175
rect 265951 293147 265999 293175
rect 265689 293113 265999 293147
rect 265689 293085 265737 293113
rect 265765 293085 265799 293113
rect 265827 293085 265861 293113
rect 265889 293085 265923 293113
rect 265951 293085 265999 293113
rect 265689 293051 265999 293085
rect 265689 293023 265737 293051
rect 265765 293023 265799 293051
rect 265827 293023 265861 293051
rect 265889 293023 265923 293051
rect 265951 293023 265999 293051
rect 265689 292989 265999 293023
rect 265689 292961 265737 292989
rect 265765 292961 265799 292989
rect 265827 292961 265861 292989
rect 265889 292961 265923 292989
rect 265951 292961 265999 292989
rect 265689 284175 265999 292961
rect 275926 294322 275954 294327
rect 265689 284147 265737 284175
rect 265765 284147 265799 284175
rect 265827 284147 265861 284175
rect 265889 284147 265923 284175
rect 265951 284147 265999 284175
rect 265689 284113 265999 284147
rect 265689 284085 265737 284113
rect 265765 284085 265799 284113
rect 265827 284085 265861 284113
rect 265889 284085 265923 284113
rect 265951 284085 265999 284113
rect 265689 284051 265999 284085
rect 265689 284023 265737 284051
rect 265765 284023 265799 284051
rect 265827 284023 265861 284051
rect 265889 284023 265923 284051
rect 265951 284023 265999 284051
rect 265689 283989 265999 284023
rect 265689 283961 265737 283989
rect 265765 283961 265799 283989
rect 265827 283961 265861 283989
rect 265889 283961 265923 283989
rect 265951 283961 265999 283989
rect 265689 275175 265999 283961
rect 265689 275147 265737 275175
rect 265765 275147 265799 275175
rect 265827 275147 265861 275175
rect 265889 275147 265923 275175
rect 265951 275147 265999 275175
rect 265689 275113 265999 275147
rect 265689 275085 265737 275113
rect 265765 275085 265799 275113
rect 265827 275085 265861 275113
rect 265889 275085 265923 275113
rect 265951 275085 265999 275113
rect 265689 275051 265999 275085
rect 265689 275023 265737 275051
rect 265765 275023 265799 275051
rect 265827 275023 265861 275051
rect 265889 275023 265923 275051
rect 265951 275023 265999 275051
rect 265689 274989 265999 275023
rect 265689 274961 265737 274989
rect 265765 274961 265799 274989
rect 265827 274961 265861 274989
rect 265889 274961 265923 274989
rect 265951 274961 265999 274989
rect 265689 266175 265999 274961
rect 265689 266147 265737 266175
rect 265765 266147 265799 266175
rect 265827 266147 265861 266175
rect 265889 266147 265923 266175
rect 265951 266147 265999 266175
rect 265689 266113 265999 266147
rect 265689 266085 265737 266113
rect 265765 266085 265799 266113
rect 265827 266085 265861 266113
rect 265889 266085 265923 266113
rect 265951 266085 265999 266113
rect 265689 266051 265999 266085
rect 265689 266023 265737 266051
rect 265765 266023 265799 266051
rect 265827 266023 265861 266051
rect 265889 266023 265923 266051
rect 265951 266023 265999 266051
rect 265689 265989 265999 266023
rect 265689 265961 265737 265989
rect 265765 265961 265799 265989
rect 265827 265961 265861 265989
rect 265889 265961 265923 265989
rect 265951 265961 265999 265989
rect 265689 257175 265999 265961
rect 265689 257147 265737 257175
rect 265765 257147 265799 257175
rect 265827 257147 265861 257175
rect 265889 257147 265923 257175
rect 265951 257147 265999 257175
rect 265689 257113 265999 257147
rect 265689 257085 265737 257113
rect 265765 257085 265799 257113
rect 265827 257085 265861 257113
rect 265889 257085 265923 257113
rect 265951 257085 265999 257113
rect 265689 257051 265999 257085
rect 265689 257023 265737 257051
rect 265765 257023 265799 257051
rect 265827 257023 265861 257051
rect 265889 257023 265923 257051
rect 265951 257023 265999 257051
rect 265689 256989 265999 257023
rect 265689 256961 265737 256989
rect 265765 256961 265799 256989
rect 265827 256961 265861 256989
rect 265889 256961 265923 256989
rect 265951 256961 265999 256989
rect 265689 248175 265999 256961
rect 265689 248147 265737 248175
rect 265765 248147 265799 248175
rect 265827 248147 265861 248175
rect 265889 248147 265923 248175
rect 265951 248147 265999 248175
rect 265689 248113 265999 248147
rect 265689 248085 265737 248113
rect 265765 248085 265799 248113
rect 265827 248085 265861 248113
rect 265889 248085 265923 248113
rect 265951 248085 265999 248113
rect 265689 248051 265999 248085
rect 265689 248023 265737 248051
rect 265765 248023 265799 248051
rect 265827 248023 265861 248051
rect 265889 248023 265923 248051
rect 265951 248023 265999 248051
rect 265689 247989 265999 248023
rect 265689 247961 265737 247989
rect 265765 247961 265799 247989
rect 265827 247961 265861 247989
rect 265889 247961 265923 247989
rect 265951 247961 265999 247989
rect 265689 239175 265999 247961
rect 265689 239147 265737 239175
rect 265765 239147 265799 239175
rect 265827 239147 265861 239175
rect 265889 239147 265923 239175
rect 265951 239147 265999 239175
rect 265689 239113 265999 239147
rect 265689 239085 265737 239113
rect 265765 239085 265799 239113
rect 265827 239085 265861 239113
rect 265889 239085 265923 239113
rect 265951 239085 265999 239113
rect 265689 239051 265999 239085
rect 265689 239023 265737 239051
rect 265765 239023 265799 239051
rect 265827 239023 265861 239051
rect 265889 239023 265923 239051
rect 265951 239023 265999 239051
rect 265689 238989 265999 239023
rect 265689 238961 265737 238989
rect 265765 238961 265799 238989
rect 265827 238961 265861 238989
rect 265889 238961 265923 238989
rect 265951 238961 265999 238989
rect 265689 230175 265999 238961
rect 265689 230147 265737 230175
rect 265765 230147 265799 230175
rect 265827 230147 265861 230175
rect 265889 230147 265923 230175
rect 265951 230147 265999 230175
rect 265689 230113 265999 230147
rect 265689 230085 265737 230113
rect 265765 230085 265799 230113
rect 265827 230085 265861 230113
rect 265889 230085 265923 230113
rect 265951 230085 265999 230113
rect 265689 230051 265999 230085
rect 265689 230023 265737 230051
rect 265765 230023 265799 230051
rect 265827 230023 265861 230051
rect 265889 230023 265923 230051
rect 265951 230023 265999 230051
rect 265689 229989 265999 230023
rect 265689 229961 265737 229989
rect 265765 229961 265799 229989
rect 265827 229961 265861 229989
rect 265889 229961 265923 229989
rect 265951 229961 265999 229989
rect 265689 221175 265999 229961
rect 265689 221147 265737 221175
rect 265765 221147 265799 221175
rect 265827 221147 265861 221175
rect 265889 221147 265923 221175
rect 265951 221147 265999 221175
rect 265689 221113 265999 221147
rect 265689 221085 265737 221113
rect 265765 221085 265799 221113
rect 265827 221085 265861 221113
rect 265889 221085 265923 221113
rect 265951 221085 265999 221113
rect 265689 221051 265999 221085
rect 265689 221023 265737 221051
rect 265765 221023 265799 221051
rect 265827 221023 265861 221051
rect 265889 221023 265923 221051
rect 265951 221023 265999 221051
rect 265689 220989 265999 221023
rect 265689 220961 265737 220989
rect 265765 220961 265799 220989
rect 265827 220961 265861 220989
rect 265889 220961 265923 220989
rect 265951 220961 265999 220989
rect 265689 212175 265999 220961
rect 265689 212147 265737 212175
rect 265765 212147 265799 212175
rect 265827 212147 265861 212175
rect 265889 212147 265923 212175
rect 265951 212147 265999 212175
rect 265689 212113 265999 212147
rect 265689 212085 265737 212113
rect 265765 212085 265799 212113
rect 265827 212085 265861 212113
rect 265889 212085 265923 212113
rect 265951 212085 265999 212113
rect 265689 212051 265999 212085
rect 265689 212023 265737 212051
rect 265765 212023 265799 212051
rect 265827 212023 265861 212051
rect 265889 212023 265923 212051
rect 265951 212023 265999 212051
rect 265689 211989 265999 212023
rect 265689 211961 265737 211989
rect 265765 211961 265799 211989
rect 265827 211961 265861 211989
rect 265889 211961 265923 211989
rect 265951 211961 265999 211989
rect 265689 203175 265999 211961
rect 265689 203147 265737 203175
rect 265765 203147 265799 203175
rect 265827 203147 265861 203175
rect 265889 203147 265923 203175
rect 265951 203147 265999 203175
rect 265689 203113 265999 203147
rect 265689 203085 265737 203113
rect 265765 203085 265799 203113
rect 265827 203085 265861 203113
rect 265889 203085 265923 203113
rect 265951 203085 265999 203113
rect 265689 203051 265999 203085
rect 265689 203023 265737 203051
rect 265765 203023 265799 203051
rect 265827 203023 265861 203051
rect 265889 203023 265923 203051
rect 265951 203023 265999 203051
rect 265689 202989 265999 203023
rect 265689 202961 265737 202989
rect 265765 202961 265799 202989
rect 265827 202961 265861 202989
rect 265889 202961 265923 202989
rect 265951 202961 265999 202989
rect 265689 194175 265999 202961
rect 265689 194147 265737 194175
rect 265765 194147 265799 194175
rect 265827 194147 265861 194175
rect 265889 194147 265923 194175
rect 265951 194147 265999 194175
rect 265689 194113 265999 194147
rect 265689 194085 265737 194113
rect 265765 194085 265799 194113
rect 265827 194085 265861 194113
rect 265889 194085 265923 194113
rect 265951 194085 265999 194113
rect 265689 194051 265999 194085
rect 265689 194023 265737 194051
rect 265765 194023 265799 194051
rect 265827 194023 265861 194051
rect 265889 194023 265923 194051
rect 265951 194023 265999 194051
rect 265689 193989 265999 194023
rect 265689 193961 265737 193989
rect 265765 193961 265799 193989
rect 265827 193961 265861 193989
rect 265889 193961 265923 193989
rect 265951 193961 265999 193989
rect 265689 185175 265999 193961
rect 265689 185147 265737 185175
rect 265765 185147 265799 185175
rect 265827 185147 265861 185175
rect 265889 185147 265923 185175
rect 265951 185147 265999 185175
rect 265689 185113 265999 185147
rect 265689 185085 265737 185113
rect 265765 185085 265799 185113
rect 265827 185085 265861 185113
rect 265889 185085 265923 185113
rect 265951 185085 265999 185113
rect 265689 185051 265999 185085
rect 265689 185023 265737 185051
rect 265765 185023 265799 185051
rect 265827 185023 265861 185051
rect 265889 185023 265923 185051
rect 265951 185023 265999 185051
rect 265689 184989 265999 185023
rect 265689 184961 265737 184989
rect 265765 184961 265799 184989
rect 265827 184961 265861 184989
rect 265889 184961 265923 184989
rect 265951 184961 265999 184989
rect 265689 176175 265999 184961
rect 265689 176147 265737 176175
rect 265765 176147 265799 176175
rect 265827 176147 265861 176175
rect 265889 176147 265923 176175
rect 265951 176147 265999 176175
rect 265689 176113 265999 176147
rect 265689 176085 265737 176113
rect 265765 176085 265799 176113
rect 265827 176085 265861 176113
rect 265889 176085 265923 176113
rect 265951 176085 265999 176113
rect 265689 176051 265999 176085
rect 265689 176023 265737 176051
rect 265765 176023 265799 176051
rect 265827 176023 265861 176051
rect 265889 176023 265923 176051
rect 265951 176023 265999 176051
rect 265689 175989 265999 176023
rect 265689 175961 265737 175989
rect 265765 175961 265799 175989
rect 265827 175961 265861 175989
rect 265889 175961 265923 175989
rect 265951 175961 265999 175989
rect 265689 167175 265999 175961
rect 265689 167147 265737 167175
rect 265765 167147 265799 167175
rect 265827 167147 265861 167175
rect 265889 167147 265923 167175
rect 265951 167147 265999 167175
rect 265689 167113 265999 167147
rect 265689 167085 265737 167113
rect 265765 167085 265799 167113
rect 265827 167085 265861 167113
rect 265889 167085 265923 167113
rect 265951 167085 265999 167113
rect 265689 167051 265999 167085
rect 265689 167023 265737 167051
rect 265765 167023 265799 167051
rect 265827 167023 265861 167051
rect 265889 167023 265923 167051
rect 265951 167023 265999 167051
rect 265689 166989 265999 167023
rect 265689 166961 265737 166989
rect 265765 166961 265799 166989
rect 265827 166961 265861 166989
rect 265889 166961 265923 166989
rect 265951 166961 265999 166989
rect 265689 158175 265999 166961
rect 265689 158147 265737 158175
rect 265765 158147 265799 158175
rect 265827 158147 265861 158175
rect 265889 158147 265923 158175
rect 265951 158147 265999 158175
rect 265689 158113 265999 158147
rect 265689 158085 265737 158113
rect 265765 158085 265799 158113
rect 265827 158085 265861 158113
rect 265889 158085 265923 158113
rect 265951 158085 265999 158113
rect 265689 158051 265999 158085
rect 265689 158023 265737 158051
rect 265765 158023 265799 158051
rect 265827 158023 265861 158051
rect 265889 158023 265923 158051
rect 265951 158023 265999 158051
rect 265689 157989 265999 158023
rect 265689 157961 265737 157989
rect 265765 157961 265799 157989
rect 265827 157961 265861 157989
rect 265889 157961 265923 157989
rect 265951 157961 265999 157989
rect 265689 149175 265999 157961
rect 271726 287714 271754 287719
rect 271726 157234 271754 287686
rect 275086 274498 275114 274503
rect 272566 254674 272594 254679
rect 271726 157201 271754 157206
rect 271782 208418 271810 208423
rect 265689 149147 265737 149175
rect 265765 149147 265799 149175
rect 265827 149147 265861 149175
rect 265889 149147 265923 149175
rect 265951 149147 265999 149175
rect 265689 149113 265999 149147
rect 265689 149085 265737 149113
rect 265765 149085 265799 149113
rect 265827 149085 265861 149113
rect 265889 149085 265923 149113
rect 265951 149085 265999 149113
rect 265689 149051 265999 149085
rect 265689 149023 265737 149051
rect 265765 149023 265799 149051
rect 265827 149023 265861 149051
rect 265889 149023 265923 149051
rect 265951 149023 265999 149051
rect 265689 148989 265999 149023
rect 265689 148961 265737 148989
rect 265765 148961 265799 148989
rect 265827 148961 265861 148989
rect 265889 148961 265923 148989
rect 265951 148961 265999 148989
rect 265689 140175 265999 148961
rect 271726 155554 271754 155559
rect 271726 148274 271754 155526
rect 271782 151858 271810 208390
rect 271782 151825 271810 151830
rect 271838 188594 271866 188599
rect 271838 150514 271866 188566
rect 271838 150481 271866 150486
rect 271894 175378 271922 175383
rect 271894 149618 271922 175350
rect 271894 149585 271922 149590
rect 271950 168770 271978 168775
rect 271950 149170 271978 168742
rect 272566 154994 272594 254646
rect 272566 154961 272594 154966
rect 272622 248066 272650 248071
rect 272622 154546 272650 248038
rect 273406 234850 273434 234855
rect 272622 154513 272650 154518
rect 272678 215082 272706 215087
rect 272678 152306 272706 215054
rect 272678 152273 272706 152278
rect 272734 181986 272762 181991
rect 272734 150066 272762 181958
rect 272734 150033 272762 150038
rect 272790 162162 272818 162167
rect 271950 149137 271978 149142
rect 272790 148722 272818 162134
rect 273406 153650 273434 234822
rect 275086 156338 275114 274470
rect 275926 157682 275954 294294
rect 279189 290175 279499 298392
rect 279189 290147 279237 290175
rect 279265 290147 279299 290175
rect 279327 290147 279361 290175
rect 279389 290147 279423 290175
rect 279451 290147 279499 290175
rect 279189 290113 279499 290147
rect 279189 290085 279237 290113
rect 279265 290085 279299 290113
rect 279327 290085 279361 290113
rect 279389 290085 279423 290113
rect 279451 290085 279499 290113
rect 279189 290051 279499 290085
rect 279189 290023 279237 290051
rect 279265 290023 279299 290051
rect 279327 290023 279361 290051
rect 279389 290023 279423 290051
rect 279451 290023 279499 290051
rect 279189 289989 279499 290023
rect 279189 289961 279237 289989
rect 279265 289961 279299 289989
rect 279327 289961 279361 289989
rect 279389 289961 279423 289989
rect 279451 289961 279499 289989
rect 279189 281175 279499 289961
rect 279189 281147 279237 281175
rect 279265 281147 279299 281175
rect 279327 281147 279361 281175
rect 279389 281147 279423 281175
rect 279451 281147 279499 281175
rect 279189 281113 279499 281147
rect 279189 281085 279237 281113
rect 279265 281085 279299 281113
rect 279327 281085 279361 281113
rect 279389 281085 279423 281113
rect 279451 281085 279499 281113
rect 279189 281051 279499 281085
rect 279189 281023 279237 281051
rect 279265 281023 279299 281051
rect 279327 281023 279361 281051
rect 279389 281023 279423 281051
rect 279451 281023 279499 281051
rect 279189 280989 279499 281023
rect 279189 280961 279237 280989
rect 279265 280961 279299 280989
rect 279327 280961 279361 280989
rect 279389 280961 279423 280989
rect 279451 280961 279499 280989
rect 279189 272175 279499 280961
rect 279189 272147 279237 272175
rect 279265 272147 279299 272175
rect 279327 272147 279361 272175
rect 279389 272147 279423 272175
rect 279451 272147 279499 272175
rect 279189 272113 279499 272147
rect 279189 272085 279237 272113
rect 279265 272085 279299 272113
rect 279327 272085 279361 272113
rect 279389 272085 279423 272113
rect 279451 272085 279499 272113
rect 279189 272051 279499 272085
rect 279189 272023 279237 272051
rect 279265 272023 279299 272051
rect 279327 272023 279361 272051
rect 279389 272023 279423 272051
rect 279451 272023 279499 272051
rect 279189 271989 279499 272023
rect 279189 271961 279237 271989
rect 279265 271961 279299 271989
rect 279327 271961 279361 271989
rect 279389 271961 279423 271989
rect 279451 271961 279499 271989
rect 278446 267890 278474 267895
rect 277606 228242 277634 228247
rect 275926 157649 275954 157654
rect 276766 195202 276794 195207
rect 275086 156305 275114 156310
rect 273406 153617 273434 153622
rect 276766 150962 276794 195174
rect 277606 153202 277634 228214
rect 278446 155890 278474 267862
rect 278446 155857 278474 155862
rect 279189 263175 279499 271961
rect 279189 263147 279237 263175
rect 279265 263147 279299 263175
rect 279327 263147 279361 263175
rect 279389 263147 279423 263175
rect 279451 263147 279499 263175
rect 279189 263113 279499 263147
rect 279189 263085 279237 263113
rect 279265 263085 279299 263113
rect 279327 263085 279361 263113
rect 279389 263085 279423 263113
rect 279451 263085 279499 263113
rect 279189 263051 279499 263085
rect 279189 263023 279237 263051
rect 279265 263023 279299 263051
rect 279327 263023 279361 263051
rect 279389 263023 279423 263051
rect 279451 263023 279499 263051
rect 279189 262989 279499 263023
rect 279189 262961 279237 262989
rect 279265 262961 279299 262989
rect 279327 262961 279361 262989
rect 279389 262961 279423 262989
rect 279451 262961 279499 262989
rect 279189 254175 279499 262961
rect 279189 254147 279237 254175
rect 279265 254147 279299 254175
rect 279327 254147 279361 254175
rect 279389 254147 279423 254175
rect 279451 254147 279499 254175
rect 279189 254113 279499 254147
rect 279189 254085 279237 254113
rect 279265 254085 279299 254113
rect 279327 254085 279361 254113
rect 279389 254085 279423 254113
rect 279451 254085 279499 254113
rect 279189 254051 279499 254085
rect 279189 254023 279237 254051
rect 279265 254023 279299 254051
rect 279327 254023 279361 254051
rect 279389 254023 279423 254051
rect 279451 254023 279499 254051
rect 279189 253989 279499 254023
rect 279189 253961 279237 253989
rect 279265 253961 279299 253989
rect 279327 253961 279361 253989
rect 279389 253961 279423 253989
rect 279451 253961 279499 253989
rect 279189 245175 279499 253961
rect 279189 245147 279237 245175
rect 279265 245147 279299 245175
rect 279327 245147 279361 245175
rect 279389 245147 279423 245175
rect 279451 245147 279499 245175
rect 279189 245113 279499 245147
rect 279189 245085 279237 245113
rect 279265 245085 279299 245113
rect 279327 245085 279361 245113
rect 279389 245085 279423 245113
rect 279451 245085 279499 245113
rect 279189 245051 279499 245085
rect 279189 245023 279237 245051
rect 279265 245023 279299 245051
rect 279327 245023 279361 245051
rect 279389 245023 279423 245051
rect 279451 245023 279499 245051
rect 279189 244989 279499 245023
rect 279189 244961 279237 244989
rect 279265 244961 279299 244989
rect 279327 244961 279361 244989
rect 279389 244961 279423 244989
rect 279451 244961 279499 244989
rect 279189 236175 279499 244961
rect 279189 236147 279237 236175
rect 279265 236147 279299 236175
rect 279327 236147 279361 236175
rect 279389 236147 279423 236175
rect 279451 236147 279499 236175
rect 279189 236113 279499 236147
rect 279189 236085 279237 236113
rect 279265 236085 279299 236113
rect 279327 236085 279361 236113
rect 279389 236085 279423 236113
rect 279451 236085 279499 236113
rect 279189 236051 279499 236085
rect 279189 236023 279237 236051
rect 279265 236023 279299 236051
rect 279327 236023 279361 236051
rect 279389 236023 279423 236051
rect 279451 236023 279499 236051
rect 279189 235989 279499 236023
rect 279189 235961 279237 235989
rect 279265 235961 279299 235989
rect 279327 235961 279361 235989
rect 279389 235961 279423 235989
rect 279451 235961 279499 235989
rect 279189 227175 279499 235961
rect 279189 227147 279237 227175
rect 279265 227147 279299 227175
rect 279327 227147 279361 227175
rect 279389 227147 279423 227175
rect 279451 227147 279499 227175
rect 279189 227113 279499 227147
rect 279189 227085 279237 227113
rect 279265 227085 279299 227113
rect 279327 227085 279361 227113
rect 279389 227085 279423 227113
rect 279451 227085 279499 227113
rect 279189 227051 279499 227085
rect 279189 227023 279237 227051
rect 279265 227023 279299 227051
rect 279327 227023 279361 227051
rect 279389 227023 279423 227051
rect 279451 227023 279499 227051
rect 279189 226989 279499 227023
rect 279189 226961 279237 226989
rect 279265 226961 279299 226989
rect 279327 226961 279361 226989
rect 279389 226961 279423 226989
rect 279451 226961 279499 226989
rect 279189 218175 279499 226961
rect 279189 218147 279237 218175
rect 279265 218147 279299 218175
rect 279327 218147 279361 218175
rect 279389 218147 279423 218175
rect 279451 218147 279499 218175
rect 279189 218113 279499 218147
rect 279189 218085 279237 218113
rect 279265 218085 279299 218113
rect 279327 218085 279361 218113
rect 279389 218085 279423 218113
rect 279451 218085 279499 218113
rect 279189 218051 279499 218085
rect 279189 218023 279237 218051
rect 279265 218023 279299 218051
rect 279327 218023 279361 218051
rect 279389 218023 279423 218051
rect 279451 218023 279499 218051
rect 279189 217989 279499 218023
rect 279189 217961 279237 217989
rect 279265 217961 279299 217989
rect 279327 217961 279361 217989
rect 279389 217961 279423 217989
rect 279451 217961 279499 217989
rect 279189 209175 279499 217961
rect 279189 209147 279237 209175
rect 279265 209147 279299 209175
rect 279327 209147 279361 209175
rect 279389 209147 279423 209175
rect 279451 209147 279499 209175
rect 279189 209113 279499 209147
rect 279189 209085 279237 209113
rect 279265 209085 279299 209113
rect 279327 209085 279361 209113
rect 279389 209085 279423 209113
rect 279451 209085 279499 209113
rect 279189 209051 279499 209085
rect 279189 209023 279237 209051
rect 279265 209023 279299 209051
rect 279327 209023 279361 209051
rect 279389 209023 279423 209051
rect 279451 209023 279499 209051
rect 279189 208989 279499 209023
rect 279189 208961 279237 208989
rect 279265 208961 279299 208989
rect 279327 208961 279361 208989
rect 279389 208961 279423 208989
rect 279451 208961 279499 208989
rect 279189 200175 279499 208961
rect 279189 200147 279237 200175
rect 279265 200147 279299 200175
rect 279327 200147 279361 200175
rect 279389 200147 279423 200175
rect 279451 200147 279499 200175
rect 279189 200113 279499 200147
rect 279189 200085 279237 200113
rect 279265 200085 279299 200113
rect 279327 200085 279361 200113
rect 279389 200085 279423 200113
rect 279451 200085 279499 200113
rect 279189 200051 279499 200085
rect 279189 200023 279237 200051
rect 279265 200023 279299 200051
rect 279327 200023 279361 200051
rect 279389 200023 279423 200051
rect 279451 200023 279499 200051
rect 279189 199989 279499 200023
rect 279189 199961 279237 199989
rect 279265 199961 279299 199989
rect 279327 199961 279361 199989
rect 279389 199961 279423 199989
rect 279451 199961 279499 199989
rect 279189 191175 279499 199961
rect 279189 191147 279237 191175
rect 279265 191147 279299 191175
rect 279327 191147 279361 191175
rect 279389 191147 279423 191175
rect 279451 191147 279499 191175
rect 279189 191113 279499 191147
rect 279189 191085 279237 191113
rect 279265 191085 279299 191113
rect 279327 191085 279361 191113
rect 279389 191085 279423 191113
rect 279451 191085 279499 191113
rect 279189 191051 279499 191085
rect 279189 191023 279237 191051
rect 279265 191023 279299 191051
rect 279327 191023 279361 191051
rect 279389 191023 279423 191051
rect 279451 191023 279499 191051
rect 279189 190989 279499 191023
rect 279189 190961 279237 190989
rect 279265 190961 279299 190989
rect 279327 190961 279361 190989
rect 279389 190961 279423 190989
rect 279451 190961 279499 190989
rect 279189 182175 279499 190961
rect 279189 182147 279237 182175
rect 279265 182147 279299 182175
rect 279327 182147 279361 182175
rect 279389 182147 279423 182175
rect 279451 182147 279499 182175
rect 279189 182113 279499 182147
rect 279189 182085 279237 182113
rect 279265 182085 279299 182113
rect 279327 182085 279361 182113
rect 279389 182085 279423 182113
rect 279451 182085 279499 182113
rect 279189 182051 279499 182085
rect 279189 182023 279237 182051
rect 279265 182023 279299 182051
rect 279327 182023 279361 182051
rect 279389 182023 279423 182051
rect 279451 182023 279499 182051
rect 279189 181989 279499 182023
rect 279189 181961 279237 181989
rect 279265 181961 279299 181989
rect 279327 181961 279361 181989
rect 279389 181961 279423 181989
rect 279451 181961 279499 181989
rect 279189 173175 279499 181961
rect 279189 173147 279237 173175
rect 279265 173147 279299 173175
rect 279327 173147 279361 173175
rect 279389 173147 279423 173175
rect 279451 173147 279499 173175
rect 279189 173113 279499 173147
rect 279189 173085 279237 173113
rect 279265 173085 279299 173113
rect 279327 173085 279361 173113
rect 279389 173085 279423 173113
rect 279451 173085 279499 173113
rect 279189 173051 279499 173085
rect 279189 173023 279237 173051
rect 279265 173023 279299 173051
rect 279327 173023 279361 173051
rect 279389 173023 279423 173051
rect 279451 173023 279499 173051
rect 279189 172989 279499 173023
rect 279189 172961 279237 172989
rect 279265 172961 279299 172989
rect 279327 172961 279361 172989
rect 279389 172961 279423 172989
rect 279451 172961 279499 172989
rect 279189 164175 279499 172961
rect 279189 164147 279237 164175
rect 279265 164147 279299 164175
rect 279327 164147 279361 164175
rect 279389 164147 279423 164175
rect 279451 164147 279499 164175
rect 279189 164113 279499 164147
rect 279189 164085 279237 164113
rect 279265 164085 279299 164113
rect 279327 164085 279361 164113
rect 279389 164085 279423 164113
rect 279451 164085 279499 164113
rect 279189 164051 279499 164085
rect 279189 164023 279237 164051
rect 279265 164023 279299 164051
rect 279327 164023 279361 164051
rect 279389 164023 279423 164051
rect 279451 164023 279499 164051
rect 279189 163989 279499 164023
rect 279189 163961 279237 163989
rect 279265 163961 279299 163989
rect 279327 163961 279361 163989
rect 279389 163961 279423 163989
rect 279451 163961 279499 163989
rect 277606 153169 277634 153174
rect 279189 155175 279499 163961
rect 279189 155147 279237 155175
rect 279265 155147 279299 155175
rect 279327 155147 279361 155175
rect 279389 155147 279423 155175
rect 279451 155147 279499 155175
rect 279189 155113 279499 155147
rect 279189 155085 279237 155113
rect 279265 155085 279299 155113
rect 279327 155085 279361 155113
rect 279389 155085 279423 155113
rect 279451 155085 279499 155113
rect 279189 155051 279499 155085
rect 279189 155023 279237 155051
rect 279265 155023 279299 155051
rect 279327 155023 279361 155051
rect 279389 155023 279423 155051
rect 279451 155023 279499 155051
rect 279189 154989 279499 155023
rect 279189 154961 279237 154989
rect 279265 154961 279299 154989
rect 279327 154961 279361 154989
rect 279389 154961 279423 154989
rect 279451 154961 279499 154989
rect 276766 150929 276794 150934
rect 272790 148689 272818 148694
rect 271726 148241 271754 148246
rect 271894 147378 271922 147383
rect 271782 146930 271810 146935
rect 265689 140147 265737 140175
rect 265765 140147 265799 140175
rect 265827 140147 265861 140175
rect 265889 140147 265923 140175
rect 265951 140147 265999 140175
rect 265689 140113 265999 140147
rect 265689 140085 265737 140113
rect 265765 140085 265799 140113
rect 265827 140085 265861 140113
rect 265889 140085 265923 140113
rect 265951 140085 265999 140113
rect 265689 140051 265999 140085
rect 265689 140023 265737 140051
rect 265765 140023 265799 140051
rect 265827 140023 265861 140051
rect 265889 140023 265923 140051
rect 265951 140023 265999 140051
rect 265689 139989 265999 140023
rect 265689 139961 265737 139989
rect 265765 139961 265799 139989
rect 265827 139961 265861 139989
rect 265889 139961 265923 139989
rect 265951 139961 265999 139989
rect 265689 131175 265999 139961
rect 265689 131147 265737 131175
rect 265765 131147 265799 131175
rect 265827 131147 265861 131175
rect 265889 131147 265923 131175
rect 265951 131147 265999 131175
rect 265689 131113 265999 131147
rect 265689 131085 265737 131113
rect 265765 131085 265799 131113
rect 265827 131085 265861 131113
rect 265889 131085 265923 131113
rect 265951 131085 265999 131113
rect 265689 131051 265999 131085
rect 265689 131023 265737 131051
rect 265765 131023 265799 131051
rect 265827 131023 265861 131051
rect 265889 131023 265923 131051
rect 265951 131023 265999 131051
rect 265689 130989 265999 131023
rect 265689 130961 265737 130989
rect 265765 130961 265799 130989
rect 265827 130961 265861 130989
rect 265889 130961 265923 130989
rect 265951 130961 265999 130989
rect 265689 125367 265999 130961
rect 271726 145586 271754 145591
rect 271726 125594 271754 145558
rect 271782 135730 271810 146902
rect 271782 135697 271810 135702
rect 271838 144242 271866 144247
rect 271838 125650 271866 144214
rect 271894 142338 271922 147350
rect 279189 146175 279499 154961
rect 279189 146147 279237 146175
rect 279265 146147 279299 146175
rect 279327 146147 279361 146175
rect 279389 146147 279423 146175
rect 279451 146147 279499 146175
rect 279189 146113 279499 146147
rect 279189 146085 279237 146113
rect 279265 146085 279299 146113
rect 279327 146085 279361 146113
rect 279389 146085 279423 146113
rect 279451 146085 279499 146113
rect 279189 146051 279499 146085
rect 276990 146034 277018 146039
rect 276934 144690 276962 144695
rect 276878 143346 276906 143351
rect 271894 142305 271922 142310
rect 271950 142898 271978 142903
rect 271950 125706 271978 142870
rect 276150 142002 276178 142007
rect 276038 140658 276066 140663
rect 275982 138866 276010 138871
rect 271950 125673 271978 125678
rect 275926 137970 275954 137975
rect 271838 125617 271866 125622
rect 271726 125561 271754 125566
rect 158169 122147 158217 122175
rect 158245 122147 158279 122175
rect 158307 122147 158341 122175
rect 158369 122147 158403 122175
rect 158431 122147 158479 122175
rect 158169 122113 158479 122147
rect 158169 122085 158217 122113
rect 158245 122085 158279 122113
rect 158307 122085 158341 122113
rect 158369 122085 158403 122113
rect 158431 122085 158479 122113
rect 158169 122051 158479 122085
rect 158169 122023 158217 122051
rect 158245 122023 158279 122051
rect 158307 122023 158341 122051
rect 158369 122023 158403 122051
rect 158431 122023 158479 122051
rect 158169 121989 158479 122023
rect 158169 121961 158217 121989
rect 158245 121961 158279 121989
rect 158307 121961 158341 121989
rect 158369 121961 158403 121989
rect 158431 121961 158479 121989
rect 158169 113175 158479 121961
rect 169904 122175 170064 122192
rect 169904 122147 169939 122175
rect 169967 122147 170001 122175
rect 170029 122147 170064 122175
rect 169904 122113 170064 122147
rect 169904 122085 169939 122113
rect 169967 122085 170001 122113
rect 170029 122085 170064 122113
rect 169904 122051 170064 122085
rect 169904 122023 169939 122051
rect 169967 122023 170001 122051
rect 170029 122023 170064 122051
rect 169904 121989 170064 122023
rect 169904 121961 169939 121989
rect 169967 121961 170001 121989
rect 170029 121961 170064 121989
rect 169904 121944 170064 121961
rect 185264 122175 185424 122192
rect 185264 122147 185299 122175
rect 185327 122147 185361 122175
rect 185389 122147 185424 122175
rect 185264 122113 185424 122147
rect 185264 122085 185299 122113
rect 185327 122085 185361 122113
rect 185389 122085 185424 122113
rect 185264 122051 185424 122085
rect 185264 122023 185299 122051
rect 185327 122023 185361 122051
rect 185389 122023 185424 122051
rect 185264 121989 185424 122023
rect 185264 121961 185299 121989
rect 185327 121961 185361 121989
rect 185389 121961 185424 121989
rect 185264 121944 185424 121961
rect 200624 122175 200784 122192
rect 200624 122147 200659 122175
rect 200687 122147 200721 122175
rect 200749 122147 200784 122175
rect 200624 122113 200784 122147
rect 200624 122085 200659 122113
rect 200687 122085 200721 122113
rect 200749 122085 200784 122113
rect 200624 122051 200784 122085
rect 200624 122023 200659 122051
rect 200687 122023 200721 122051
rect 200749 122023 200784 122051
rect 200624 121989 200784 122023
rect 200624 121961 200659 121989
rect 200687 121961 200721 121989
rect 200749 121961 200784 121989
rect 200624 121944 200784 121961
rect 215984 122175 216144 122192
rect 215984 122147 216019 122175
rect 216047 122147 216081 122175
rect 216109 122147 216144 122175
rect 215984 122113 216144 122147
rect 215984 122085 216019 122113
rect 216047 122085 216081 122113
rect 216109 122085 216144 122113
rect 215984 122051 216144 122085
rect 215984 122023 216019 122051
rect 216047 122023 216081 122051
rect 216109 122023 216144 122051
rect 215984 121989 216144 122023
rect 215984 121961 216019 121989
rect 216047 121961 216081 121989
rect 216109 121961 216144 121989
rect 215984 121944 216144 121961
rect 231344 122175 231504 122192
rect 231344 122147 231379 122175
rect 231407 122147 231441 122175
rect 231469 122147 231504 122175
rect 231344 122113 231504 122147
rect 231344 122085 231379 122113
rect 231407 122085 231441 122113
rect 231469 122085 231504 122113
rect 231344 122051 231504 122085
rect 231344 122023 231379 122051
rect 231407 122023 231441 122051
rect 231469 122023 231504 122051
rect 231344 121989 231504 122023
rect 231344 121961 231379 121989
rect 231407 121961 231441 121989
rect 231469 121961 231504 121989
rect 231344 121944 231504 121961
rect 246704 122175 246864 122192
rect 246704 122147 246739 122175
rect 246767 122147 246801 122175
rect 246829 122147 246864 122175
rect 246704 122113 246864 122147
rect 246704 122085 246739 122113
rect 246767 122085 246801 122113
rect 246829 122085 246864 122113
rect 246704 122051 246864 122085
rect 246704 122023 246739 122051
rect 246767 122023 246801 122051
rect 246829 122023 246864 122051
rect 246704 121989 246864 122023
rect 246704 121961 246739 121989
rect 246767 121961 246801 121989
rect 246829 121961 246864 121989
rect 246704 121944 246864 121961
rect 262064 122175 262224 122192
rect 262064 122147 262099 122175
rect 262127 122147 262161 122175
rect 262189 122147 262224 122175
rect 262064 122113 262224 122147
rect 262064 122085 262099 122113
rect 262127 122085 262161 122113
rect 262189 122085 262224 122113
rect 262064 122051 262224 122085
rect 262064 122023 262099 122051
rect 262127 122023 262161 122051
rect 262189 122023 262224 122051
rect 262064 121989 262224 122023
rect 262064 121961 262099 121989
rect 262127 121961 262161 121989
rect 262189 121961 262224 121989
rect 262064 121944 262224 121961
rect 162224 119175 162384 119192
rect 162224 119147 162259 119175
rect 162287 119147 162321 119175
rect 162349 119147 162384 119175
rect 162224 119113 162384 119147
rect 162224 119085 162259 119113
rect 162287 119085 162321 119113
rect 162349 119085 162384 119113
rect 162224 119051 162384 119085
rect 162224 119023 162259 119051
rect 162287 119023 162321 119051
rect 162349 119023 162384 119051
rect 162224 118989 162384 119023
rect 162224 118961 162259 118989
rect 162287 118961 162321 118989
rect 162349 118961 162384 118989
rect 162224 118944 162384 118961
rect 177584 119175 177744 119192
rect 177584 119147 177619 119175
rect 177647 119147 177681 119175
rect 177709 119147 177744 119175
rect 177584 119113 177744 119147
rect 177584 119085 177619 119113
rect 177647 119085 177681 119113
rect 177709 119085 177744 119113
rect 177584 119051 177744 119085
rect 177584 119023 177619 119051
rect 177647 119023 177681 119051
rect 177709 119023 177744 119051
rect 177584 118989 177744 119023
rect 177584 118961 177619 118989
rect 177647 118961 177681 118989
rect 177709 118961 177744 118989
rect 177584 118944 177744 118961
rect 192944 119175 193104 119192
rect 192944 119147 192979 119175
rect 193007 119147 193041 119175
rect 193069 119147 193104 119175
rect 192944 119113 193104 119147
rect 192944 119085 192979 119113
rect 193007 119085 193041 119113
rect 193069 119085 193104 119113
rect 192944 119051 193104 119085
rect 192944 119023 192979 119051
rect 193007 119023 193041 119051
rect 193069 119023 193104 119051
rect 192944 118989 193104 119023
rect 192944 118961 192979 118989
rect 193007 118961 193041 118989
rect 193069 118961 193104 118989
rect 192944 118944 193104 118961
rect 208304 119175 208464 119192
rect 208304 119147 208339 119175
rect 208367 119147 208401 119175
rect 208429 119147 208464 119175
rect 208304 119113 208464 119147
rect 208304 119085 208339 119113
rect 208367 119085 208401 119113
rect 208429 119085 208464 119113
rect 208304 119051 208464 119085
rect 208304 119023 208339 119051
rect 208367 119023 208401 119051
rect 208429 119023 208464 119051
rect 208304 118989 208464 119023
rect 208304 118961 208339 118989
rect 208367 118961 208401 118989
rect 208429 118961 208464 118989
rect 208304 118944 208464 118961
rect 223664 119175 223824 119192
rect 223664 119147 223699 119175
rect 223727 119147 223761 119175
rect 223789 119147 223824 119175
rect 223664 119113 223824 119147
rect 223664 119085 223699 119113
rect 223727 119085 223761 119113
rect 223789 119085 223824 119113
rect 223664 119051 223824 119085
rect 223664 119023 223699 119051
rect 223727 119023 223761 119051
rect 223789 119023 223824 119051
rect 223664 118989 223824 119023
rect 223664 118961 223699 118989
rect 223727 118961 223761 118989
rect 223789 118961 223824 118989
rect 223664 118944 223824 118961
rect 239024 119175 239184 119192
rect 239024 119147 239059 119175
rect 239087 119147 239121 119175
rect 239149 119147 239184 119175
rect 239024 119113 239184 119147
rect 239024 119085 239059 119113
rect 239087 119085 239121 119113
rect 239149 119085 239184 119113
rect 239024 119051 239184 119085
rect 239024 119023 239059 119051
rect 239087 119023 239121 119051
rect 239149 119023 239184 119051
rect 239024 118989 239184 119023
rect 239024 118961 239059 118989
rect 239087 118961 239121 118989
rect 239149 118961 239184 118989
rect 239024 118944 239184 118961
rect 254384 119175 254544 119192
rect 254384 119147 254419 119175
rect 254447 119147 254481 119175
rect 254509 119147 254544 119175
rect 254384 119113 254544 119147
rect 254384 119085 254419 119113
rect 254447 119085 254481 119113
rect 254509 119085 254544 119113
rect 254384 119051 254544 119085
rect 254384 119023 254419 119051
rect 254447 119023 254481 119051
rect 254509 119023 254544 119051
rect 254384 118989 254544 119023
rect 254384 118961 254419 118989
rect 254447 118961 254481 118989
rect 254509 118961 254544 118989
rect 254384 118944 254544 118961
rect 269744 119175 269904 119192
rect 269744 119147 269779 119175
rect 269807 119147 269841 119175
rect 269869 119147 269904 119175
rect 269744 119113 269904 119147
rect 269744 119085 269779 119113
rect 269807 119085 269841 119113
rect 269869 119085 269904 119113
rect 269744 119051 269904 119085
rect 269744 119023 269779 119051
rect 269807 119023 269841 119051
rect 269869 119023 269904 119051
rect 269744 118989 269904 119023
rect 269744 118961 269779 118989
rect 269807 118961 269841 118989
rect 269869 118961 269904 118989
rect 269744 118944 269904 118961
rect 158169 113147 158217 113175
rect 158245 113147 158279 113175
rect 158307 113147 158341 113175
rect 158369 113147 158403 113175
rect 158431 113147 158479 113175
rect 158169 113113 158479 113147
rect 158169 113085 158217 113113
rect 158245 113085 158279 113113
rect 158307 113085 158341 113113
rect 158369 113085 158403 113113
rect 158431 113085 158479 113113
rect 158169 113051 158479 113085
rect 158169 113023 158217 113051
rect 158245 113023 158279 113051
rect 158307 113023 158341 113051
rect 158369 113023 158403 113051
rect 158431 113023 158479 113051
rect 158169 112989 158479 113023
rect 158169 112961 158217 112989
rect 158245 112961 158279 112989
rect 158307 112961 158341 112989
rect 158369 112961 158403 112989
rect 158431 112961 158479 112989
rect 158169 104175 158479 112961
rect 169904 113175 170064 113192
rect 169904 113147 169939 113175
rect 169967 113147 170001 113175
rect 170029 113147 170064 113175
rect 169904 113113 170064 113147
rect 169904 113085 169939 113113
rect 169967 113085 170001 113113
rect 170029 113085 170064 113113
rect 169904 113051 170064 113085
rect 169904 113023 169939 113051
rect 169967 113023 170001 113051
rect 170029 113023 170064 113051
rect 169904 112989 170064 113023
rect 169904 112961 169939 112989
rect 169967 112961 170001 112989
rect 170029 112961 170064 112989
rect 169904 112944 170064 112961
rect 185264 113175 185424 113192
rect 185264 113147 185299 113175
rect 185327 113147 185361 113175
rect 185389 113147 185424 113175
rect 185264 113113 185424 113147
rect 185264 113085 185299 113113
rect 185327 113085 185361 113113
rect 185389 113085 185424 113113
rect 185264 113051 185424 113085
rect 185264 113023 185299 113051
rect 185327 113023 185361 113051
rect 185389 113023 185424 113051
rect 185264 112989 185424 113023
rect 185264 112961 185299 112989
rect 185327 112961 185361 112989
rect 185389 112961 185424 112989
rect 185264 112944 185424 112961
rect 200624 113175 200784 113192
rect 200624 113147 200659 113175
rect 200687 113147 200721 113175
rect 200749 113147 200784 113175
rect 200624 113113 200784 113147
rect 200624 113085 200659 113113
rect 200687 113085 200721 113113
rect 200749 113085 200784 113113
rect 200624 113051 200784 113085
rect 200624 113023 200659 113051
rect 200687 113023 200721 113051
rect 200749 113023 200784 113051
rect 200624 112989 200784 113023
rect 200624 112961 200659 112989
rect 200687 112961 200721 112989
rect 200749 112961 200784 112989
rect 200624 112944 200784 112961
rect 215984 113175 216144 113192
rect 215984 113147 216019 113175
rect 216047 113147 216081 113175
rect 216109 113147 216144 113175
rect 215984 113113 216144 113147
rect 215984 113085 216019 113113
rect 216047 113085 216081 113113
rect 216109 113085 216144 113113
rect 215984 113051 216144 113085
rect 215984 113023 216019 113051
rect 216047 113023 216081 113051
rect 216109 113023 216144 113051
rect 215984 112989 216144 113023
rect 215984 112961 216019 112989
rect 216047 112961 216081 112989
rect 216109 112961 216144 112989
rect 215984 112944 216144 112961
rect 231344 113175 231504 113192
rect 231344 113147 231379 113175
rect 231407 113147 231441 113175
rect 231469 113147 231504 113175
rect 231344 113113 231504 113147
rect 231344 113085 231379 113113
rect 231407 113085 231441 113113
rect 231469 113085 231504 113113
rect 231344 113051 231504 113085
rect 231344 113023 231379 113051
rect 231407 113023 231441 113051
rect 231469 113023 231504 113051
rect 231344 112989 231504 113023
rect 231344 112961 231379 112989
rect 231407 112961 231441 112989
rect 231469 112961 231504 112989
rect 231344 112944 231504 112961
rect 246704 113175 246864 113192
rect 246704 113147 246739 113175
rect 246767 113147 246801 113175
rect 246829 113147 246864 113175
rect 246704 113113 246864 113147
rect 246704 113085 246739 113113
rect 246767 113085 246801 113113
rect 246829 113085 246864 113113
rect 246704 113051 246864 113085
rect 246704 113023 246739 113051
rect 246767 113023 246801 113051
rect 246829 113023 246864 113051
rect 246704 112989 246864 113023
rect 246704 112961 246739 112989
rect 246767 112961 246801 112989
rect 246829 112961 246864 112989
rect 246704 112944 246864 112961
rect 262064 113175 262224 113192
rect 262064 113147 262099 113175
rect 262127 113147 262161 113175
rect 262189 113147 262224 113175
rect 262064 113113 262224 113147
rect 262064 113085 262099 113113
rect 262127 113085 262161 113113
rect 262189 113085 262224 113113
rect 262064 113051 262224 113085
rect 262064 113023 262099 113051
rect 262127 113023 262161 113051
rect 262189 113023 262224 113051
rect 262064 112989 262224 113023
rect 262064 112961 262099 112989
rect 262127 112961 262161 112989
rect 262189 112961 262224 112989
rect 262064 112944 262224 112961
rect 162224 110175 162384 110192
rect 162224 110147 162259 110175
rect 162287 110147 162321 110175
rect 162349 110147 162384 110175
rect 162224 110113 162384 110147
rect 162224 110085 162259 110113
rect 162287 110085 162321 110113
rect 162349 110085 162384 110113
rect 162224 110051 162384 110085
rect 162224 110023 162259 110051
rect 162287 110023 162321 110051
rect 162349 110023 162384 110051
rect 162224 109989 162384 110023
rect 162224 109961 162259 109989
rect 162287 109961 162321 109989
rect 162349 109961 162384 109989
rect 162224 109944 162384 109961
rect 177584 110175 177744 110192
rect 177584 110147 177619 110175
rect 177647 110147 177681 110175
rect 177709 110147 177744 110175
rect 177584 110113 177744 110147
rect 177584 110085 177619 110113
rect 177647 110085 177681 110113
rect 177709 110085 177744 110113
rect 177584 110051 177744 110085
rect 177584 110023 177619 110051
rect 177647 110023 177681 110051
rect 177709 110023 177744 110051
rect 177584 109989 177744 110023
rect 177584 109961 177619 109989
rect 177647 109961 177681 109989
rect 177709 109961 177744 109989
rect 177584 109944 177744 109961
rect 192944 110175 193104 110192
rect 192944 110147 192979 110175
rect 193007 110147 193041 110175
rect 193069 110147 193104 110175
rect 192944 110113 193104 110147
rect 192944 110085 192979 110113
rect 193007 110085 193041 110113
rect 193069 110085 193104 110113
rect 192944 110051 193104 110085
rect 192944 110023 192979 110051
rect 193007 110023 193041 110051
rect 193069 110023 193104 110051
rect 192944 109989 193104 110023
rect 192944 109961 192979 109989
rect 193007 109961 193041 109989
rect 193069 109961 193104 109989
rect 192944 109944 193104 109961
rect 208304 110175 208464 110192
rect 208304 110147 208339 110175
rect 208367 110147 208401 110175
rect 208429 110147 208464 110175
rect 208304 110113 208464 110147
rect 208304 110085 208339 110113
rect 208367 110085 208401 110113
rect 208429 110085 208464 110113
rect 208304 110051 208464 110085
rect 208304 110023 208339 110051
rect 208367 110023 208401 110051
rect 208429 110023 208464 110051
rect 208304 109989 208464 110023
rect 208304 109961 208339 109989
rect 208367 109961 208401 109989
rect 208429 109961 208464 109989
rect 208304 109944 208464 109961
rect 223664 110175 223824 110192
rect 223664 110147 223699 110175
rect 223727 110147 223761 110175
rect 223789 110147 223824 110175
rect 223664 110113 223824 110147
rect 223664 110085 223699 110113
rect 223727 110085 223761 110113
rect 223789 110085 223824 110113
rect 223664 110051 223824 110085
rect 223664 110023 223699 110051
rect 223727 110023 223761 110051
rect 223789 110023 223824 110051
rect 223664 109989 223824 110023
rect 223664 109961 223699 109989
rect 223727 109961 223761 109989
rect 223789 109961 223824 109989
rect 223664 109944 223824 109961
rect 239024 110175 239184 110192
rect 239024 110147 239059 110175
rect 239087 110147 239121 110175
rect 239149 110147 239184 110175
rect 239024 110113 239184 110147
rect 239024 110085 239059 110113
rect 239087 110085 239121 110113
rect 239149 110085 239184 110113
rect 239024 110051 239184 110085
rect 239024 110023 239059 110051
rect 239087 110023 239121 110051
rect 239149 110023 239184 110051
rect 239024 109989 239184 110023
rect 239024 109961 239059 109989
rect 239087 109961 239121 109989
rect 239149 109961 239184 109989
rect 239024 109944 239184 109961
rect 254384 110175 254544 110192
rect 254384 110147 254419 110175
rect 254447 110147 254481 110175
rect 254509 110147 254544 110175
rect 254384 110113 254544 110147
rect 254384 110085 254419 110113
rect 254447 110085 254481 110113
rect 254509 110085 254544 110113
rect 254384 110051 254544 110085
rect 254384 110023 254419 110051
rect 254447 110023 254481 110051
rect 254509 110023 254544 110051
rect 254384 109989 254544 110023
rect 254384 109961 254419 109989
rect 254447 109961 254481 109989
rect 254509 109961 254544 109989
rect 254384 109944 254544 109961
rect 269744 110175 269904 110192
rect 269744 110147 269779 110175
rect 269807 110147 269841 110175
rect 269869 110147 269904 110175
rect 269744 110113 269904 110147
rect 269744 110085 269779 110113
rect 269807 110085 269841 110113
rect 269869 110085 269904 110113
rect 269744 110051 269904 110085
rect 269744 110023 269779 110051
rect 269807 110023 269841 110051
rect 269869 110023 269904 110051
rect 269744 109989 269904 110023
rect 269744 109961 269779 109989
rect 269807 109961 269841 109989
rect 269869 109961 269904 109989
rect 269744 109944 269904 109961
rect 158169 104147 158217 104175
rect 158245 104147 158279 104175
rect 158307 104147 158341 104175
rect 158369 104147 158403 104175
rect 158431 104147 158479 104175
rect 158169 104113 158479 104147
rect 158169 104085 158217 104113
rect 158245 104085 158279 104113
rect 158307 104085 158341 104113
rect 158369 104085 158403 104113
rect 158431 104085 158479 104113
rect 158169 104051 158479 104085
rect 158169 104023 158217 104051
rect 158245 104023 158279 104051
rect 158307 104023 158341 104051
rect 158369 104023 158403 104051
rect 158431 104023 158479 104051
rect 158169 103989 158479 104023
rect 158169 103961 158217 103989
rect 158245 103961 158279 103989
rect 158307 103961 158341 103989
rect 158369 103961 158403 103989
rect 158431 103961 158479 103989
rect 158169 95175 158479 103961
rect 169904 104175 170064 104192
rect 169904 104147 169939 104175
rect 169967 104147 170001 104175
rect 170029 104147 170064 104175
rect 169904 104113 170064 104147
rect 169904 104085 169939 104113
rect 169967 104085 170001 104113
rect 170029 104085 170064 104113
rect 169904 104051 170064 104085
rect 169904 104023 169939 104051
rect 169967 104023 170001 104051
rect 170029 104023 170064 104051
rect 169904 103989 170064 104023
rect 169904 103961 169939 103989
rect 169967 103961 170001 103989
rect 170029 103961 170064 103989
rect 169904 103944 170064 103961
rect 185264 104175 185424 104192
rect 185264 104147 185299 104175
rect 185327 104147 185361 104175
rect 185389 104147 185424 104175
rect 185264 104113 185424 104147
rect 185264 104085 185299 104113
rect 185327 104085 185361 104113
rect 185389 104085 185424 104113
rect 185264 104051 185424 104085
rect 185264 104023 185299 104051
rect 185327 104023 185361 104051
rect 185389 104023 185424 104051
rect 185264 103989 185424 104023
rect 185264 103961 185299 103989
rect 185327 103961 185361 103989
rect 185389 103961 185424 103989
rect 185264 103944 185424 103961
rect 200624 104175 200784 104192
rect 200624 104147 200659 104175
rect 200687 104147 200721 104175
rect 200749 104147 200784 104175
rect 200624 104113 200784 104147
rect 200624 104085 200659 104113
rect 200687 104085 200721 104113
rect 200749 104085 200784 104113
rect 200624 104051 200784 104085
rect 200624 104023 200659 104051
rect 200687 104023 200721 104051
rect 200749 104023 200784 104051
rect 200624 103989 200784 104023
rect 200624 103961 200659 103989
rect 200687 103961 200721 103989
rect 200749 103961 200784 103989
rect 200624 103944 200784 103961
rect 215984 104175 216144 104192
rect 215984 104147 216019 104175
rect 216047 104147 216081 104175
rect 216109 104147 216144 104175
rect 215984 104113 216144 104147
rect 215984 104085 216019 104113
rect 216047 104085 216081 104113
rect 216109 104085 216144 104113
rect 215984 104051 216144 104085
rect 215984 104023 216019 104051
rect 216047 104023 216081 104051
rect 216109 104023 216144 104051
rect 215984 103989 216144 104023
rect 215984 103961 216019 103989
rect 216047 103961 216081 103989
rect 216109 103961 216144 103989
rect 215984 103944 216144 103961
rect 231344 104175 231504 104192
rect 231344 104147 231379 104175
rect 231407 104147 231441 104175
rect 231469 104147 231504 104175
rect 231344 104113 231504 104147
rect 231344 104085 231379 104113
rect 231407 104085 231441 104113
rect 231469 104085 231504 104113
rect 231344 104051 231504 104085
rect 231344 104023 231379 104051
rect 231407 104023 231441 104051
rect 231469 104023 231504 104051
rect 231344 103989 231504 104023
rect 231344 103961 231379 103989
rect 231407 103961 231441 103989
rect 231469 103961 231504 103989
rect 231344 103944 231504 103961
rect 246704 104175 246864 104192
rect 246704 104147 246739 104175
rect 246767 104147 246801 104175
rect 246829 104147 246864 104175
rect 246704 104113 246864 104147
rect 246704 104085 246739 104113
rect 246767 104085 246801 104113
rect 246829 104085 246864 104113
rect 246704 104051 246864 104085
rect 246704 104023 246739 104051
rect 246767 104023 246801 104051
rect 246829 104023 246864 104051
rect 246704 103989 246864 104023
rect 246704 103961 246739 103989
rect 246767 103961 246801 103989
rect 246829 103961 246864 103989
rect 246704 103944 246864 103961
rect 262064 104175 262224 104192
rect 262064 104147 262099 104175
rect 262127 104147 262161 104175
rect 262189 104147 262224 104175
rect 262064 104113 262224 104147
rect 262064 104085 262099 104113
rect 262127 104085 262161 104113
rect 262189 104085 262224 104113
rect 262064 104051 262224 104085
rect 262064 104023 262099 104051
rect 262127 104023 262161 104051
rect 262189 104023 262224 104051
rect 262064 103989 262224 104023
rect 262064 103961 262099 103989
rect 262127 103961 262161 103989
rect 262189 103961 262224 103989
rect 262064 103944 262224 103961
rect 162224 101175 162384 101192
rect 162224 101147 162259 101175
rect 162287 101147 162321 101175
rect 162349 101147 162384 101175
rect 162224 101113 162384 101147
rect 162224 101085 162259 101113
rect 162287 101085 162321 101113
rect 162349 101085 162384 101113
rect 162224 101051 162384 101085
rect 162224 101023 162259 101051
rect 162287 101023 162321 101051
rect 162349 101023 162384 101051
rect 162224 100989 162384 101023
rect 162224 100961 162259 100989
rect 162287 100961 162321 100989
rect 162349 100961 162384 100989
rect 162224 100944 162384 100961
rect 177584 101175 177744 101192
rect 177584 101147 177619 101175
rect 177647 101147 177681 101175
rect 177709 101147 177744 101175
rect 177584 101113 177744 101147
rect 177584 101085 177619 101113
rect 177647 101085 177681 101113
rect 177709 101085 177744 101113
rect 177584 101051 177744 101085
rect 177584 101023 177619 101051
rect 177647 101023 177681 101051
rect 177709 101023 177744 101051
rect 177584 100989 177744 101023
rect 177584 100961 177619 100989
rect 177647 100961 177681 100989
rect 177709 100961 177744 100989
rect 177584 100944 177744 100961
rect 192944 101175 193104 101192
rect 192944 101147 192979 101175
rect 193007 101147 193041 101175
rect 193069 101147 193104 101175
rect 192944 101113 193104 101147
rect 192944 101085 192979 101113
rect 193007 101085 193041 101113
rect 193069 101085 193104 101113
rect 192944 101051 193104 101085
rect 192944 101023 192979 101051
rect 193007 101023 193041 101051
rect 193069 101023 193104 101051
rect 192944 100989 193104 101023
rect 192944 100961 192979 100989
rect 193007 100961 193041 100989
rect 193069 100961 193104 100989
rect 192944 100944 193104 100961
rect 208304 101175 208464 101192
rect 208304 101147 208339 101175
rect 208367 101147 208401 101175
rect 208429 101147 208464 101175
rect 208304 101113 208464 101147
rect 208304 101085 208339 101113
rect 208367 101085 208401 101113
rect 208429 101085 208464 101113
rect 208304 101051 208464 101085
rect 208304 101023 208339 101051
rect 208367 101023 208401 101051
rect 208429 101023 208464 101051
rect 208304 100989 208464 101023
rect 208304 100961 208339 100989
rect 208367 100961 208401 100989
rect 208429 100961 208464 100989
rect 208304 100944 208464 100961
rect 223664 101175 223824 101192
rect 223664 101147 223699 101175
rect 223727 101147 223761 101175
rect 223789 101147 223824 101175
rect 223664 101113 223824 101147
rect 223664 101085 223699 101113
rect 223727 101085 223761 101113
rect 223789 101085 223824 101113
rect 223664 101051 223824 101085
rect 223664 101023 223699 101051
rect 223727 101023 223761 101051
rect 223789 101023 223824 101051
rect 223664 100989 223824 101023
rect 223664 100961 223699 100989
rect 223727 100961 223761 100989
rect 223789 100961 223824 100989
rect 223664 100944 223824 100961
rect 239024 101175 239184 101192
rect 239024 101147 239059 101175
rect 239087 101147 239121 101175
rect 239149 101147 239184 101175
rect 239024 101113 239184 101147
rect 239024 101085 239059 101113
rect 239087 101085 239121 101113
rect 239149 101085 239184 101113
rect 239024 101051 239184 101085
rect 239024 101023 239059 101051
rect 239087 101023 239121 101051
rect 239149 101023 239184 101051
rect 239024 100989 239184 101023
rect 239024 100961 239059 100989
rect 239087 100961 239121 100989
rect 239149 100961 239184 100989
rect 239024 100944 239184 100961
rect 254384 101175 254544 101192
rect 254384 101147 254419 101175
rect 254447 101147 254481 101175
rect 254509 101147 254544 101175
rect 254384 101113 254544 101147
rect 254384 101085 254419 101113
rect 254447 101085 254481 101113
rect 254509 101085 254544 101113
rect 254384 101051 254544 101085
rect 254384 101023 254419 101051
rect 254447 101023 254481 101051
rect 254509 101023 254544 101051
rect 254384 100989 254544 101023
rect 254384 100961 254419 100989
rect 254447 100961 254481 100989
rect 254509 100961 254544 100989
rect 254384 100944 254544 100961
rect 269744 101175 269904 101192
rect 269744 101147 269779 101175
rect 269807 101147 269841 101175
rect 269869 101147 269904 101175
rect 269744 101113 269904 101147
rect 269744 101085 269779 101113
rect 269807 101085 269841 101113
rect 269869 101085 269904 101113
rect 269744 101051 269904 101085
rect 269744 101023 269779 101051
rect 269807 101023 269841 101051
rect 269869 101023 269904 101051
rect 269744 100989 269904 101023
rect 269744 100961 269779 100989
rect 269807 100961 269841 100989
rect 269869 100961 269904 100989
rect 269744 100944 269904 100961
rect 158169 95147 158217 95175
rect 158245 95147 158279 95175
rect 158307 95147 158341 95175
rect 158369 95147 158403 95175
rect 158431 95147 158479 95175
rect 158169 95113 158479 95147
rect 158169 95085 158217 95113
rect 158245 95085 158279 95113
rect 158307 95085 158341 95113
rect 158369 95085 158403 95113
rect 158431 95085 158479 95113
rect 158169 95051 158479 95085
rect 158169 95023 158217 95051
rect 158245 95023 158279 95051
rect 158307 95023 158341 95051
rect 158369 95023 158403 95051
rect 158431 95023 158479 95051
rect 158169 94989 158479 95023
rect 158169 94961 158217 94989
rect 158245 94961 158279 94989
rect 158307 94961 158341 94989
rect 158369 94961 158403 94989
rect 158431 94961 158479 94989
rect 158169 86175 158479 94961
rect 169904 95175 170064 95192
rect 169904 95147 169939 95175
rect 169967 95147 170001 95175
rect 170029 95147 170064 95175
rect 169904 95113 170064 95147
rect 169904 95085 169939 95113
rect 169967 95085 170001 95113
rect 170029 95085 170064 95113
rect 169904 95051 170064 95085
rect 169904 95023 169939 95051
rect 169967 95023 170001 95051
rect 170029 95023 170064 95051
rect 169904 94989 170064 95023
rect 169904 94961 169939 94989
rect 169967 94961 170001 94989
rect 170029 94961 170064 94989
rect 169904 94944 170064 94961
rect 185264 95175 185424 95192
rect 185264 95147 185299 95175
rect 185327 95147 185361 95175
rect 185389 95147 185424 95175
rect 185264 95113 185424 95147
rect 185264 95085 185299 95113
rect 185327 95085 185361 95113
rect 185389 95085 185424 95113
rect 185264 95051 185424 95085
rect 185264 95023 185299 95051
rect 185327 95023 185361 95051
rect 185389 95023 185424 95051
rect 185264 94989 185424 95023
rect 185264 94961 185299 94989
rect 185327 94961 185361 94989
rect 185389 94961 185424 94989
rect 185264 94944 185424 94961
rect 200624 95175 200784 95192
rect 200624 95147 200659 95175
rect 200687 95147 200721 95175
rect 200749 95147 200784 95175
rect 200624 95113 200784 95147
rect 200624 95085 200659 95113
rect 200687 95085 200721 95113
rect 200749 95085 200784 95113
rect 200624 95051 200784 95085
rect 200624 95023 200659 95051
rect 200687 95023 200721 95051
rect 200749 95023 200784 95051
rect 200624 94989 200784 95023
rect 200624 94961 200659 94989
rect 200687 94961 200721 94989
rect 200749 94961 200784 94989
rect 200624 94944 200784 94961
rect 215984 95175 216144 95192
rect 215984 95147 216019 95175
rect 216047 95147 216081 95175
rect 216109 95147 216144 95175
rect 215984 95113 216144 95147
rect 215984 95085 216019 95113
rect 216047 95085 216081 95113
rect 216109 95085 216144 95113
rect 215984 95051 216144 95085
rect 215984 95023 216019 95051
rect 216047 95023 216081 95051
rect 216109 95023 216144 95051
rect 215984 94989 216144 95023
rect 215984 94961 216019 94989
rect 216047 94961 216081 94989
rect 216109 94961 216144 94989
rect 215984 94944 216144 94961
rect 231344 95175 231504 95192
rect 231344 95147 231379 95175
rect 231407 95147 231441 95175
rect 231469 95147 231504 95175
rect 231344 95113 231504 95147
rect 231344 95085 231379 95113
rect 231407 95085 231441 95113
rect 231469 95085 231504 95113
rect 231344 95051 231504 95085
rect 231344 95023 231379 95051
rect 231407 95023 231441 95051
rect 231469 95023 231504 95051
rect 231344 94989 231504 95023
rect 231344 94961 231379 94989
rect 231407 94961 231441 94989
rect 231469 94961 231504 94989
rect 231344 94944 231504 94961
rect 246704 95175 246864 95192
rect 246704 95147 246739 95175
rect 246767 95147 246801 95175
rect 246829 95147 246864 95175
rect 246704 95113 246864 95147
rect 246704 95085 246739 95113
rect 246767 95085 246801 95113
rect 246829 95085 246864 95113
rect 246704 95051 246864 95085
rect 246704 95023 246739 95051
rect 246767 95023 246801 95051
rect 246829 95023 246864 95051
rect 246704 94989 246864 95023
rect 246704 94961 246739 94989
rect 246767 94961 246801 94989
rect 246829 94961 246864 94989
rect 246704 94944 246864 94961
rect 262064 95175 262224 95192
rect 262064 95147 262099 95175
rect 262127 95147 262161 95175
rect 262189 95147 262224 95175
rect 262064 95113 262224 95147
rect 262064 95085 262099 95113
rect 262127 95085 262161 95113
rect 262189 95085 262224 95113
rect 262064 95051 262224 95085
rect 262064 95023 262099 95051
rect 262127 95023 262161 95051
rect 262189 95023 262224 95051
rect 262064 94989 262224 95023
rect 262064 94961 262099 94989
rect 262127 94961 262161 94989
rect 262189 94961 262224 94989
rect 262064 94944 262224 94961
rect 162224 92175 162384 92192
rect 162224 92147 162259 92175
rect 162287 92147 162321 92175
rect 162349 92147 162384 92175
rect 162224 92113 162384 92147
rect 162224 92085 162259 92113
rect 162287 92085 162321 92113
rect 162349 92085 162384 92113
rect 162224 92051 162384 92085
rect 162224 92023 162259 92051
rect 162287 92023 162321 92051
rect 162349 92023 162384 92051
rect 162224 91989 162384 92023
rect 162224 91961 162259 91989
rect 162287 91961 162321 91989
rect 162349 91961 162384 91989
rect 162224 91944 162384 91961
rect 177584 92175 177744 92192
rect 177584 92147 177619 92175
rect 177647 92147 177681 92175
rect 177709 92147 177744 92175
rect 177584 92113 177744 92147
rect 177584 92085 177619 92113
rect 177647 92085 177681 92113
rect 177709 92085 177744 92113
rect 177584 92051 177744 92085
rect 177584 92023 177619 92051
rect 177647 92023 177681 92051
rect 177709 92023 177744 92051
rect 177584 91989 177744 92023
rect 177584 91961 177619 91989
rect 177647 91961 177681 91989
rect 177709 91961 177744 91989
rect 177584 91944 177744 91961
rect 192944 92175 193104 92192
rect 192944 92147 192979 92175
rect 193007 92147 193041 92175
rect 193069 92147 193104 92175
rect 192944 92113 193104 92147
rect 192944 92085 192979 92113
rect 193007 92085 193041 92113
rect 193069 92085 193104 92113
rect 192944 92051 193104 92085
rect 192944 92023 192979 92051
rect 193007 92023 193041 92051
rect 193069 92023 193104 92051
rect 192944 91989 193104 92023
rect 192944 91961 192979 91989
rect 193007 91961 193041 91989
rect 193069 91961 193104 91989
rect 192944 91944 193104 91961
rect 208304 92175 208464 92192
rect 208304 92147 208339 92175
rect 208367 92147 208401 92175
rect 208429 92147 208464 92175
rect 208304 92113 208464 92147
rect 208304 92085 208339 92113
rect 208367 92085 208401 92113
rect 208429 92085 208464 92113
rect 208304 92051 208464 92085
rect 208304 92023 208339 92051
rect 208367 92023 208401 92051
rect 208429 92023 208464 92051
rect 208304 91989 208464 92023
rect 208304 91961 208339 91989
rect 208367 91961 208401 91989
rect 208429 91961 208464 91989
rect 208304 91944 208464 91961
rect 223664 92175 223824 92192
rect 223664 92147 223699 92175
rect 223727 92147 223761 92175
rect 223789 92147 223824 92175
rect 223664 92113 223824 92147
rect 223664 92085 223699 92113
rect 223727 92085 223761 92113
rect 223789 92085 223824 92113
rect 223664 92051 223824 92085
rect 223664 92023 223699 92051
rect 223727 92023 223761 92051
rect 223789 92023 223824 92051
rect 223664 91989 223824 92023
rect 223664 91961 223699 91989
rect 223727 91961 223761 91989
rect 223789 91961 223824 91989
rect 223664 91944 223824 91961
rect 239024 92175 239184 92192
rect 239024 92147 239059 92175
rect 239087 92147 239121 92175
rect 239149 92147 239184 92175
rect 239024 92113 239184 92147
rect 239024 92085 239059 92113
rect 239087 92085 239121 92113
rect 239149 92085 239184 92113
rect 239024 92051 239184 92085
rect 239024 92023 239059 92051
rect 239087 92023 239121 92051
rect 239149 92023 239184 92051
rect 239024 91989 239184 92023
rect 239024 91961 239059 91989
rect 239087 91961 239121 91989
rect 239149 91961 239184 91989
rect 239024 91944 239184 91961
rect 254384 92175 254544 92192
rect 254384 92147 254419 92175
rect 254447 92147 254481 92175
rect 254509 92147 254544 92175
rect 254384 92113 254544 92147
rect 254384 92085 254419 92113
rect 254447 92085 254481 92113
rect 254509 92085 254544 92113
rect 254384 92051 254544 92085
rect 254384 92023 254419 92051
rect 254447 92023 254481 92051
rect 254509 92023 254544 92051
rect 254384 91989 254544 92023
rect 254384 91961 254419 91989
rect 254447 91961 254481 91989
rect 254509 91961 254544 91989
rect 254384 91944 254544 91961
rect 269744 92175 269904 92192
rect 269744 92147 269779 92175
rect 269807 92147 269841 92175
rect 269869 92147 269904 92175
rect 269744 92113 269904 92147
rect 269744 92085 269779 92113
rect 269807 92085 269841 92113
rect 269869 92085 269904 92113
rect 269744 92051 269904 92085
rect 269744 92023 269779 92051
rect 269807 92023 269841 92051
rect 269869 92023 269904 92051
rect 269744 91989 269904 92023
rect 269744 91961 269779 91989
rect 269807 91961 269841 91989
rect 269869 91961 269904 91989
rect 269744 91944 269904 91961
rect 158169 86147 158217 86175
rect 158245 86147 158279 86175
rect 158307 86147 158341 86175
rect 158369 86147 158403 86175
rect 158431 86147 158479 86175
rect 158169 86113 158479 86147
rect 158169 86085 158217 86113
rect 158245 86085 158279 86113
rect 158307 86085 158341 86113
rect 158369 86085 158403 86113
rect 158431 86085 158479 86113
rect 158169 86051 158479 86085
rect 158169 86023 158217 86051
rect 158245 86023 158279 86051
rect 158307 86023 158341 86051
rect 158369 86023 158403 86051
rect 158431 86023 158479 86051
rect 158169 85989 158479 86023
rect 158169 85961 158217 85989
rect 158245 85961 158279 85989
rect 158307 85961 158341 85989
rect 158369 85961 158403 85989
rect 158431 85961 158479 85989
rect 158169 77175 158479 85961
rect 169904 86175 170064 86192
rect 169904 86147 169939 86175
rect 169967 86147 170001 86175
rect 170029 86147 170064 86175
rect 169904 86113 170064 86147
rect 169904 86085 169939 86113
rect 169967 86085 170001 86113
rect 170029 86085 170064 86113
rect 169904 86051 170064 86085
rect 169904 86023 169939 86051
rect 169967 86023 170001 86051
rect 170029 86023 170064 86051
rect 169904 85989 170064 86023
rect 169904 85961 169939 85989
rect 169967 85961 170001 85989
rect 170029 85961 170064 85989
rect 169904 85944 170064 85961
rect 185264 86175 185424 86192
rect 185264 86147 185299 86175
rect 185327 86147 185361 86175
rect 185389 86147 185424 86175
rect 185264 86113 185424 86147
rect 185264 86085 185299 86113
rect 185327 86085 185361 86113
rect 185389 86085 185424 86113
rect 185264 86051 185424 86085
rect 185264 86023 185299 86051
rect 185327 86023 185361 86051
rect 185389 86023 185424 86051
rect 185264 85989 185424 86023
rect 185264 85961 185299 85989
rect 185327 85961 185361 85989
rect 185389 85961 185424 85989
rect 185264 85944 185424 85961
rect 200624 86175 200784 86192
rect 200624 86147 200659 86175
rect 200687 86147 200721 86175
rect 200749 86147 200784 86175
rect 200624 86113 200784 86147
rect 200624 86085 200659 86113
rect 200687 86085 200721 86113
rect 200749 86085 200784 86113
rect 200624 86051 200784 86085
rect 200624 86023 200659 86051
rect 200687 86023 200721 86051
rect 200749 86023 200784 86051
rect 200624 85989 200784 86023
rect 200624 85961 200659 85989
rect 200687 85961 200721 85989
rect 200749 85961 200784 85989
rect 200624 85944 200784 85961
rect 215984 86175 216144 86192
rect 215984 86147 216019 86175
rect 216047 86147 216081 86175
rect 216109 86147 216144 86175
rect 215984 86113 216144 86147
rect 215984 86085 216019 86113
rect 216047 86085 216081 86113
rect 216109 86085 216144 86113
rect 215984 86051 216144 86085
rect 215984 86023 216019 86051
rect 216047 86023 216081 86051
rect 216109 86023 216144 86051
rect 215984 85989 216144 86023
rect 215984 85961 216019 85989
rect 216047 85961 216081 85989
rect 216109 85961 216144 85989
rect 215984 85944 216144 85961
rect 231344 86175 231504 86192
rect 231344 86147 231379 86175
rect 231407 86147 231441 86175
rect 231469 86147 231504 86175
rect 231344 86113 231504 86147
rect 231344 86085 231379 86113
rect 231407 86085 231441 86113
rect 231469 86085 231504 86113
rect 231344 86051 231504 86085
rect 231344 86023 231379 86051
rect 231407 86023 231441 86051
rect 231469 86023 231504 86051
rect 231344 85989 231504 86023
rect 231344 85961 231379 85989
rect 231407 85961 231441 85989
rect 231469 85961 231504 85989
rect 231344 85944 231504 85961
rect 246704 86175 246864 86192
rect 246704 86147 246739 86175
rect 246767 86147 246801 86175
rect 246829 86147 246864 86175
rect 246704 86113 246864 86147
rect 246704 86085 246739 86113
rect 246767 86085 246801 86113
rect 246829 86085 246864 86113
rect 246704 86051 246864 86085
rect 246704 86023 246739 86051
rect 246767 86023 246801 86051
rect 246829 86023 246864 86051
rect 246704 85989 246864 86023
rect 246704 85961 246739 85989
rect 246767 85961 246801 85989
rect 246829 85961 246864 85989
rect 246704 85944 246864 85961
rect 262064 86175 262224 86192
rect 262064 86147 262099 86175
rect 262127 86147 262161 86175
rect 262189 86147 262224 86175
rect 262064 86113 262224 86147
rect 262064 86085 262099 86113
rect 262127 86085 262161 86113
rect 262189 86085 262224 86113
rect 262064 86051 262224 86085
rect 262064 86023 262099 86051
rect 262127 86023 262161 86051
rect 262189 86023 262224 86051
rect 262064 85989 262224 86023
rect 262064 85961 262099 85989
rect 262127 85961 262161 85989
rect 262189 85961 262224 85989
rect 262064 85944 262224 85961
rect 162224 83175 162384 83192
rect 162224 83147 162259 83175
rect 162287 83147 162321 83175
rect 162349 83147 162384 83175
rect 162224 83113 162384 83147
rect 162224 83085 162259 83113
rect 162287 83085 162321 83113
rect 162349 83085 162384 83113
rect 162224 83051 162384 83085
rect 162224 83023 162259 83051
rect 162287 83023 162321 83051
rect 162349 83023 162384 83051
rect 162224 82989 162384 83023
rect 162224 82961 162259 82989
rect 162287 82961 162321 82989
rect 162349 82961 162384 82989
rect 162224 82944 162384 82961
rect 177584 83175 177744 83192
rect 177584 83147 177619 83175
rect 177647 83147 177681 83175
rect 177709 83147 177744 83175
rect 177584 83113 177744 83147
rect 177584 83085 177619 83113
rect 177647 83085 177681 83113
rect 177709 83085 177744 83113
rect 177584 83051 177744 83085
rect 177584 83023 177619 83051
rect 177647 83023 177681 83051
rect 177709 83023 177744 83051
rect 177584 82989 177744 83023
rect 177584 82961 177619 82989
rect 177647 82961 177681 82989
rect 177709 82961 177744 82989
rect 177584 82944 177744 82961
rect 192944 83175 193104 83192
rect 192944 83147 192979 83175
rect 193007 83147 193041 83175
rect 193069 83147 193104 83175
rect 192944 83113 193104 83147
rect 192944 83085 192979 83113
rect 193007 83085 193041 83113
rect 193069 83085 193104 83113
rect 192944 83051 193104 83085
rect 192944 83023 192979 83051
rect 193007 83023 193041 83051
rect 193069 83023 193104 83051
rect 192944 82989 193104 83023
rect 192944 82961 192979 82989
rect 193007 82961 193041 82989
rect 193069 82961 193104 82989
rect 192944 82944 193104 82961
rect 208304 83175 208464 83192
rect 208304 83147 208339 83175
rect 208367 83147 208401 83175
rect 208429 83147 208464 83175
rect 208304 83113 208464 83147
rect 208304 83085 208339 83113
rect 208367 83085 208401 83113
rect 208429 83085 208464 83113
rect 208304 83051 208464 83085
rect 208304 83023 208339 83051
rect 208367 83023 208401 83051
rect 208429 83023 208464 83051
rect 208304 82989 208464 83023
rect 208304 82961 208339 82989
rect 208367 82961 208401 82989
rect 208429 82961 208464 82989
rect 208304 82944 208464 82961
rect 223664 83175 223824 83192
rect 223664 83147 223699 83175
rect 223727 83147 223761 83175
rect 223789 83147 223824 83175
rect 223664 83113 223824 83147
rect 223664 83085 223699 83113
rect 223727 83085 223761 83113
rect 223789 83085 223824 83113
rect 223664 83051 223824 83085
rect 223664 83023 223699 83051
rect 223727 83023 223761 83051
rect 223789 83023 223824 83051
rect 223664 82989 223824 83023
rect 223664 82961 223699 82989
rect 223727 82961 223761 82989
rect 223789 82961 223824 82989
rect 223664 82944 223824 82961
rect 239024 83175 239184 83192
rect 239024 83147 239059 83175
rect 239087 83147 239121 83175
rect 239149 83147 239184 83175
rect 239024 83113 239184 83147
rect 239024 83085 239059 83113
rect 239087 83085 239121 83113
rect 239149 83085 239184 83113
rect 239024 83051 239184 83085
rect 239024 83023 239059 83051
rect 239087 83023 239121 83051
rect 239149 83023 239184 83051
rect 239024 82989 239184 83023
rect 239024 82961 239059 82989
rect 239087 82961 239121 82989
rect 239149 82961 239184 82989
rect 239024 82944 239184 82961
rect 254384 83175 254544 83192
rect 254384 83147 254419 83175
rect 254447 83147 254481 83175
rect 254509 83147 254544 83175
rect 254384 83113 254544 83147
rect 254384 83085 254419 83113
rect 254447 83085 254481 83113
rect 254509 83085 254544 83113
rect 254384 83051 254544 83085
rect 254384 83023 254419 83051
rect 254447 83023 254481 83051
rect 254509 83023 254544 83051
rect 254384 82989 254544 83023
rect 254384 82961 254419 82989
rect 254447 82961 254481 82989
rect 254509 82961 254544 82989
rect 254384 82944 254544 82961
rect 269744 83175 269904 83192
rect 269744 83147 269779 83175
rect 269807 83147 269841 83175
rect 269869 83147 269904 83175
rect 269744 83113 269904 83147
rect 269744 83085 269779 83113
rect 269807 83085 269841 83113
rect 269869 83085 269904 83113
rect 269744 83051 269904 83085
rect 269744 83023 269779 83051
rect 269807 83023 269841 83051
rect 269869 83023 269904 83051
rect 269744 82989 269904 83023
rect 269744 82961 269779 82989
rect 269807 82961 269841 82989
rect 269869 82961 269904 82989
rect 269744 82944 269904 82961
rect 158169 77147 158217 77175
rect 158245 77147 158279 77175
rect 158307 77147 158341 77175
rect 158369 77147 158403 77175
rect 158431 77147 158479 77175
rect 158169 77113 158479 77147
rect 158169 77085 158217 77113
rect 158245 77085 158279 77113
rect 158307 77085 158341 77113
rect 158369 77085 158403 77113
rect 158431 77085 158479 77113
rect 158169 77051 158479 77085
rect 158169 77023 158217 77051
rect 158245 77023 158279 77051
rect 158307 77023 158341 77051
rect 158369 77023 158403 77051
rect 158431 77023 158479 77051
rect 158169 76989 158479 77023
rect 158169 76961 158217 76989
rect 158245 76961 158279 76989
rect 158307 76961 158341 76989
rect 158369 76961 158403 76989
rect 158431 76961 158479 76989
rect 158169 68175 158479 76961
rect 169904 77175 170064 77192
rect 169904 77147 169939 77175
rect 169967 77147 170001 77175
rect 170029 77147 170064 77175
rect 169904 77113 170064 77147
rect 169904 77085 169939 77113
rect 169967 77085 170001 77113
rect 170029 77085 170064 77113
rect 169904 77051 170064 77085
rect 169904 77023 169939 77051
rect 169967 77023 170001 77051
rect 170029 77023 170064 77051
rect 169904 76989 170064 77023
rect 169904 76961 169939 76989
rect 169967 76961 170001 76989
rect 170029 76961 170064 76989
rect 169904 76944 170064 76961
rect 185264 77175 185424 77192
rect 185264 77147 185299 77175
rect 185327 77147 185361 77175
rect 185389 77147 185424 77175
rect 185264 77113 185424 77147
rect 185264 77085 185299 77113
rect 185327 77085 185361 77113
rect 185389 77085 185424 77113
rect 185264 77051 185424 77085
rect 185264 77023 185299 77051
rect 185327 77023 185361 77051
rect 185389 77023 185424 77051
rect 185264 76989 185424 77023
rect 185264 76961 185299 76989
rect 185327 76961 185361 76989
rect 185389 76961 185424 76989
rect 185264 76944 185424 76961
rect 200624 77175 200784 77192
rect 200624 77147 200659 77175
rect 200687 77147 200721 77175
rect 200749 77147 200784 77175
rect 200624 77113 200784 77147
rect 200624 77085 200659 77113
rect 200687 77085 200721 77113
rect 200749 77085 200784 77113
rect 200624 77051 200784 77085
rect 200624 77023 200659 77051
rect 200687 77023 200721 77051
rect 200749 77023 200784 77051
rect 200624 76989 200784 77023
rect 200624 76961 200659 76989
rect 200687 76961 200721 76989
rect 200749 76961 200784 76989
rect 200624 76944 200784 76961
rect 215984 77175 216144 77192
rect 215984 77147 216019 77175
rect 216047 77147 216081 77175
rect 216109 77147 216144 77175
rect 215984 77113 216144 77147
rect 215984 77085 216019 77113
rect 216047 77085 216081 77113
rect 216109 77085 216144 77113
rect 215984 77051 216144 77085
rect 215984 77023 216019 77051
rect 216047 77023 216081 77051
rect 216109 77023 216144 77051
rect 215984 76989 216144 77023
rect 215984 76961 216019 76989
rect 216047 76961 216081 76989
rect 216109 76961 216144 76989
rect 215984 76944 216144 76961
rect 231344 77175 231504 77192
rect 231344 77147 231379 77175
rect 231407 77147 231441 77175
rect 231469 77147 231504 77175
rect 231344 77113 231504 77147
rect 231344 77085 231379 77113
rect 231407 77085 231441 77113
rect 231469 77085 231504 77113
rect 231344 77051 231504 77085
rect 231344 77023 231379 77051
rect 231407 77023 231441 77051
rect 231469 77023 231504 77051
rect 231344 76989 231504 77023
rect 231344 76961 231379 76989
rect 231407 76961 231441 76989
rect 231469 76961 231504 76989
rect 231344 76944 231504 76961
rect 246704 77175 246864 77192
rect 246704 77147 246739 77175
rect 246767 77147 246801 77175
rect 246829 77147 246864 77175
rect 246704 77113 246864 77147
rect 246704 77085 246739 77113
rect 246767 77085 246801 77113
rect 246829 77085 246864 77113
rect 246704 77051 246864 77085
rect 246704 77023 246739 77051
rect 246767 77023 246801 77051
rect 246829 77023 246864 77051
rect 246704 76989 246864 77023
rect 246704 76961 246739 76989
rect 246767 76961 246801 76989
rect 246829 76961 246864 76989
rect 246704 76944 246864 76961
rect 262064 77175 262224 77192
rect 262064 77147 262099 77175
rect 262127 77147 262161 77175
rect 262189 77147 262224 77175
rect 262064 77113 262224 77147
rect 262064 77085 262099 77113
rect 262127 77085 262161 77113
rect 262189 77085 262224 77113
rect 262064 77051 262224 77085
rect 262064 77023 262099 77051
rect 262127 77023 262161 77051
rect 262189 77023 262224 77051
rect 262064 76989 262224 77023
rect 262064 76961 262099 76989
rect 262127 76961 262161 76989
rect 262189 76961 262224 76989
rect 262064 76944 262224 76961
rect 162224 74175 162384 74192
rect 162224 74147 162259 74175
rect 162287 74147 162321 74175
rect 162349 74147 162384 74175
rect 162224 74113 162384 74147
rect 162224 74085 162259 74113
rect 162287 74085 162321 74113
rect 162349 74085 162384 74113
rect 162224 74051 162384 74085
rect 162224 74023 162259 74051
rect 162287 74023 162321 74051
rect 162349 74023 162384 74051
rect 162224 73989 162384 74023
rect 162224 73961 162259 73989
rect 162287 73961 162321 73989
rect 162349 73961 162384 73989
rect 162224 73944 162384 73961
rect 177584 74175 177744 74192
rect 177584 74147 177619 74175
rect 177647 74147 177681 74175
rect 177709 74147 177744 74175
rect 177584 74113 177744 74147
rect 177584 74085 177619 74113
rect 177647 74085 177681 74113
rect 177709 74085 177744 74113
rect 177584 74051 177744 74085
rect 177584 74023 177619 74051
rect 177647 74023 177681 74051
rect 177709 74023 177744 74051
rect 177584 73989 177744 74023
rect 177584 73961 177619 73989
rect 177647 73961 177681 73989
rect 177709 73961 177744 73989
rect 177584 73944 177744 73961
rect 192944 74175 193104 74192
rect 192944 74147 192979 74175
rect 193007 74147 193041 74175
rect 193069 74147 193104 74175
rect 192944 74113 193104 74147
rect 192944 74085 192979 74113
rect 193007 74085 193041 74113
rect 193069 74085 193104 74113
rect 192944 74051 193104 74085
rect 192944 74023 192979 74051
rect 193007 74023 193041 74051
rect 193069 74023 193104 74051
rect 192944 73989 193104 74023
rect 192944 73961 192979 73989
rect 193007 73961 193041 73989
rect 193069 73961 193104 73989
rect 192944 73944 193104 73961
rect 208304 74175 208464 74192
rect 208304 74147 208339 74175
rect 208367 74147 208401 74175
rect 208429 74147 208464 74175
rect 208304 74113 208464 74147
rect 208304 74085 208339 74113
rect 208367 74085 208401 74113
rect 208429 74085 208464 74113
rect 208304 74051 208464 74085
rect 208304 74023 208339 74051
rect 208367 74023 208401 74051
rect 208429 74023 208464 74051
rect 208304 73989 208464 74023
rect 208304 73961 208339 73989
rect 208367 73961 208401 73989
rect 208429 73961 208464 73989
rect 208304 73944 208464 73961
rect 223664 74175 223824 74192
rect 223664 74147 223699 74175
rect 223727 74147 223761 74175
rect 223789 74147 223824 74175
rect 223664 74113 223824 74147
rect 223664 74085 223699 74113
rect 223727 74085 223761 74113
rect 223789 74085 223824 74113
rect 223664 74051 223824 74085
rect 223664 74023 223699 74051
rect 223727 74023 223761 74051
rect 223789 74023 223824 74051
rect 223664 73989 223824 74023
rect 223664 73961 223699 73989
rect 223727 73961 223761 73989
rect 223789 73961 223824 73989
rect 223664 73944 223824 73961
rect 239024 74175 239184 74192
rect 239024 74147 239059 74175
rect 239087 74147 239121 74175
rect 239149 74147 239184 74175
rect 239024 74113 239184 74147
rect 239024 74085 239059 74113
rect 239087 74085 239121 74113
rect 239149 74085 239184 74113
rect 239024 74051 239184 74085
rect 239024 74023 239059 74051
rect 239087 74023 239121 74051
rect 239149 74023 239184 74051
rect 239024 73989 239184 74023
rect 239024 73961 239059 73989
rect 239087 73961 239121 73989
rect 239149 73961 239184 73989
rect 239024 73944 239184 73961
rect 254384 74175 254544 74192
rect 254384 74147 254419 74175
rect 254447 74147 254481 74175
rect 254509 74147 254544 74175
rect 254384 74113 254544 74147
rect 254384 74085 254419 74113
rect 254447 74085 254481 74113
rect 254509 74085 254544 74113
rect 254384 74051 254544 74085
rect 254384 74023 254419 74051
rect 254447 74023 254481 74051
rect 254509 74023 254544 74051
rect 254384 73989 254544 74023
rect 254384 73961 254419 73989
rect 254447 73961 254481 73989
rect 254509 73961 254544 73989
rect 254384 73944 254544 73961
rect 269744 74175 269904 74192
rect 269744 74147 269779 74175
rect 269807 74147 269841 74175
rect 269869 74147 269904 74175
rect 269744 74113 269904 74147
rect 269744 74085 269779 74113
rect 269807 74085 269841 74113
rect 269869 74085 269904 74113
rect 269744 74051 269904 74085
rect 269744 74023 269779 74051
rect 269807 74023 269841 74051
rect 269869 74023 269904 74051
rect 269744 73989 269904 74023
rect 269744 73961 269779 73989
rect 269807 73961 269841 73989
rect 269869 73961 269904 73989
rect 269744 73944 269904 73961
rect 158169 68147 158217 68175
rect 158245 68147 158279 68175
rect 158307 68147 158341 68175
rect 158369 68147 158403 68175
rect 158431 68147 158479 68175
rect 158169 68113 158479 68147
rect 158169 68085 158217 68113
rect 158245 68085 158279 68113
rect 158307 68085 158341 68113
rect 158369 68085 158403 68113
rect 158431 68085 158479 68113
rect 158169 68051 158479 68085
rect 158169 68023 158217 68051
rect 158245 68023 158279 68051
rect 158307 68023 158341 68051
rect 158369 68023 158403 68051
rect 158431 68023 158479 68051
rect 158169 67989 158479 68023
rect 158169 67961 158217 67989
rect 158245 67961 158279 67989
rect 158307 67961 158341 67989
rect 158369 67961 158403 67989
rect 158431 67961 158479 67989
rect 158169 59175 158479 67961
rect 169904 68175 170064 68192
rect 169904 68147 169939 68175
rect 169967 68147 170001 68175
rect 170029 68147 170064 68175
rect 169904 68113 170064 68147
rect 169904 68085 169939 68113
rect 169967 68085 170001 68113
rect 170029 68085 170064 68113
rect 169904 68051 170064 68085
rect 169904 68023 169939 68051
rect 169967 68023 170001 68051
rect 170029 68023 170064 68051
rect 169904 67989 170064 68023
rect 169904 67961 169939 67989
rect 169967 67961 170001 67989
rect 170029 67961 170064 67989
rect 169904 67944 170064 67961
rect 185264 68175 185424 68192
rect 185264 68147 185299 68175
rect 185327 68147 185361 68175
rect 185389 68147 185424 68175
rect 185264 68113 185424 68147
rect 185264 68085 185299 68113
rect 185327 68085 185361 68113
rect 185389 68085 185424 68113
rect 185264 68051 185424 68085
rect 185264 68023 185299 68051
rect 185327 68023 185361 68051
rect 185389 68023 185424 68051
rect 185264 67989 185424 68023
rect 185264 67961 185299 67989
rect 185327 67961 185361 67989
rect 185389 67961 185424 67989
rect 185264 67944 185424 67961
rect 200624 68175 200784 68192
rect 200624 68147 200659 68175
rect 200687 68147 200721 68175
rect 200749 68147 200784 68175
rect 200624 68113 200784 68147
rect 200624 68085 200659 68113
rect 200687 68085 200721 68113
rect 200749 68085 200784 68113
rect 200624 68051 200784 68085
rect 200624 68023 200659 68051
rect 200687 68023 200721 68051
rect 200749 68023 200784 68051
rect 200624 67989 200784 68023
rect 200624 67961 200659 67989
rect 200687 67961 200721 67989
rect 200749 67961 200784 67989
rect 200624 67944 200784 67961
rect 215984 68175 216144 68192
rect 215984 68147 216019 68175
rect 216047 68147 216081 68175
rect 216109 68147 216144 68175
rect 215984 68113 216144 68147
rect 215984 68085 216019 68113
rect 216047 68085 216081 68113
rect 216109 68085 216144 68113
rect 215984 68051 216144 68085
rect 215984 68023 216019 68051
rect 216047 68023 216081 68051
rect 216109 68023 216144 68051
rect 215984 67989 216144 68023
rect 215984 67961 216019 67989
rect 216047 67961 216081 67989
rect 216109 67961 216144 67989
rect 215984 67944 216144 67961
rect 231344 68175 231504 68192
rect 231344 68147 231379 68175
rect 231407 68147 231441 68175
rect 231469 68147 231504 68175
rect 231344 68113 231504 68147
rect 231344 68085 231379 68113
rect 231407 68085 231441 68113
rect 231469 68085 231504 68113
rect 231344 68051 231504 68085
rect 231344 68023 231379 68051
rect 231407 68023 231441 68051
rect 231469 68023 231504 68051
rect 231344 67989 231504 68023
rect 231344 67961 231379 67989
rect 231407 67961 231441 67989
rect 231469 67961 231504 67989
rect 231344 67944 231504 67961
rect 246704 68175 246864 68192
rect 246704 68147 246739 68175
rect 246767 68147 246801 68175
rect 246829 68147 246864 68175
rect 246704 68113 246864 68147
rect 246704 68085 246739 68113
rect 246767 68085 246801 68113
rect 246829 68085 246864 68113
rect 246704 68051 246864 68085
rect 246704 68023 246739 68051
rect 246767 68023 246801 68051
rect 246829 68023 246864 68051
rect 246704 67989 246864 68023
rect 246704 67961 246739 67989
rect 246767 67961 246801 67989
rect 246829 67961 246864 67989
rect 246704 67944 246864 67961
rect 262064 68175 262224 68192
rect 262064 68147 262099 68175
rect 262127 68147 262161 68175
rect 262189 68147 262224 68175
rect 262064 68113 262224 68147
rect 262064 68085 262099 68113
rect 262127 68085 262161 68113
rect 262189 68085 262224 68113
rect 262064 68051 262224 68085
rect 262064 68023 262099 68051
rect 262127 68023 262161 68051
rect 262189 68023 262224 68051
rect 262064 67989 262224 68023
rect 262064 67961 262099 67989
rect 262127 67961 262161 67989
rect 262189 67961 262224 67989
rect 262064 67944 262224 67961
rect 162224 65175 162384 65192
rect 162224 65147 162259 65175
rect 162287 65147 162321 65175
rect 162349 65147 162384 65175
rect 162224 65113 162384 65147
rect 162224 65085 162259 65113
rect 162287 65085 162321 65113
rect 162349 65085 162384 65113
rect 162224 65051 162384 65085
rect 162224 65023 162259 65051
rect 162287 65023 162321 65051
rect 162349 65023 162384 65051
rect 162224 64989 162384 65023
rect 162224 64961 162259 64989
rect 162287 64961 162321 64989
rect 162349 64961 162384 64989
rect 162224 64944 162384 64961
rect 177584 65175 177744 65192
rect 177584 65147 177619 65175
rect 177647 65147 177681 65175
rect 177709 65147 177744 65175
rect 177584 65113 177744 65147
rect 177584 65085 177619 65113
rect 177647 65085 177681 65113
rect 177709 65085 177744 65113
rect 177584 65051 177744 65085
rect 177584 65023 177619 65051
rect 177647 65023 177681 65051
rect 177709 65023 177744 65051
rect 177584 64989 177744 65023
rect 177584 64961 177619 64989
rect 177647 64961 177681 64989
rect 177709 64961 177744 64989
rect 177584 64944 177744 64961
rect 192944 65175 193104 65192
rect 192944 65147 192979 65175
rect 193007 65147 193041 65175
rect 193069 65147 193104 65175
rect 192944 65113 193104 65147
rect 192944 65085 192979 65113
rect 193007 65085 193041 65113
rect 193069 65085 193104 65113
rect 192944 65051 193104 65085
rect 192944 65023 192979 65051
rect 193007 65023 193041 65051
rect 193069 65023 193104 65051
rect 192944 64989 193104 65023
rect 192944 64961 192979 64989
rect 193007 64961 193041 64989
rect 193069 64961 193104 64989
rect 192944 64944 193104 64961
rect 208304 65175 208464 65192
rect 208304 65147 208339 65175
rect 208367 65147 208401 65175
rect 208429 65147 208464 65175
rect 208304 65113 208464 65147
rect 208304 65085 208339 65113
rect 208367 65085 208401 65113
rect 208429 65085 208464 65113
rect 208304 65051 208464 65085
rect 208304 65023 208339 65051
rect 208367 65023 208401 65051
rect 208429 65023 208464 65051
rect 208304 64989 208464 65023
rect 208304 64961 208339 64989
rect 208367 64961 208401 64989
rect 208429 64961 208464 64989
rect 208304 64944 208464 64961
rect 223664 65175 223824 65192
rect 223664 65147 223699 65175
rect 223727 65147 223761 65175
rect 223789 65147 223824 65175
rect 223664 65113 223824 65147
rect 223664 65085 223699 65113
rect 223727 65085 223761 65113
rect 223789 65085 223824 65113
rect 223664 65051 223824 65085
rect 223664 65023 223699 65051
rect 223727 65023 223761 65051
rect 223789 65023 223824 65051
rect 223664 64989 223824 65023
rect 223664 64961 223699 64989
rect 223727 64961 223761 64989
rect 223789 64961 223824 64989
rect 223664 64944 223824 64961
rect 239024 65175 239184 65192
rect 239024 65147 239059 65175
rect 239087 65147 239121 65175
rect 239149 65147 239184 65175
rect 239024 65113 239184 65147
rect 239024 65085 239059 65113
rect 239087 65085 239121 65113
rect 239149 65085 239184 65113
rect 239024 65051 239184 65085
rect 239024 65023 239059 65051
rect 239087 65023 239121 65051
rect 239149 65023 239184 65051
rect 239024 64989 239184 65023
rect 239024 64961 239059 64989
rect 239087 64961 239121 64989
rect 239149 64961 239184 64989
rect 239024 64944 239184 64961
rect 254384 65175 254544 65192
rect 254384 65147 254419 65175
rect 254447 65147 254481 65175
rect 254509 65147 254544 65175
rect 254384 65113 254544 65147
rect 254384 65085 254419 65113
rect 254447 65085 254481 65113
rect 254509 65085 254544 65113
rect 254384 65051 254544 65085
rect 254384 65023 254419 65051
rect 254447 65023 254481 65051
rect 254509 65023 254544 65051
rect 254384 64989 254544 65023
rect 254384 64961 254419 64989
rect 254447 64961 254481 64989
rect 254509 64961 254544 64989
rect 254384 64944 254544 64961
rect 269744 65175 269904 65192
rect 269744 65147 269779 65175
rect 269807 65147 269841 65175
rect 269869 65147 269904 65175
rect 269744 65113 269904 65147
rect 269744 65085 269779 65113
rect 269807 65085 269841 65113
rect 269869 65085 269904 65113
rect 269744 65051 269904 65085
rect 269744 65023 269779 65051
rect 269807 65023 269841 65051
rect 269869 65023 269904 65051
rect 269744 64989 269904 65023
rect 269744 64961 269779 64989
rect 269807 64961 269841 64989
rect 269869 64961 269904 64989
rect 269744 64944 269904 64961
rect 158169 59147 158217 59175
rect 158245 59147 158279 59175
rect 158307 59147 158341 59175
rect 158369 59147 158403 59175
rect 158431 59147 158479 59175
rect 158169 59113 158479 59147
rect 158169 59085 158217 59113
rect 158245 59085 158279 59113
rect 158307 59085 158341 59113
rect 158369 59085 158403 59113
rect 158431 59085 158479 59113
rect 158169 59051 158479 59085
rect 158169 59023 158217 59051
rect 158245 59023 158279 59051
rect 158307 59023 158341 59051
rect 158369 59023 158403 59051
rect 158431 59023 158479 59051
rect 158169 58989 158479 59023
rect 158169 58961 158217 58989
rect 158245 58961 158279 58989
rect 158307 58961 158341 58989
rect 158369 58961 158403 58989
rect 158431 58961 158479 58989
rect 158169 50175 158479 58961
rect 169904 59175 170064 59192
rect 169904 59147 169939 59175
rect 169967 59147 170001 59175
rect 170029 59147 170064 59175
rect 169904 59113 170064 59147
rect 169904 59085 169939 59113
rect 169967 59085 170001 59113
rect 170029 59085 170064 59113
rect 169904 59051 170064 59085
rect 169904 59023 169939 59051
rect 169967 59023 170001 59051
rect 170029 59023 170064 59051
rect 169904 58989 170064 59023
rect 169904 58961 169939 58989
rect 169967 58961 170001 58989
rect 170029 58961 170064 58989
rect 169904 58944 170064 58961
rect 185264 59175 185424 59192
rect 185264 59147 185299 59175
rect 185327 59147 185361 59175
rect 185389 59147 185424 59175
rect 185264 59113 185424 59147
rect 185264 59085 185299 59113
rect 185327 59085 185361 59113
rect 185389 59085 185424 59113
rect 185264 59051 185424 59085
rect 185264 59023 185299 59051
rect 185327 59023 185361 59051
rect 185389 59023 185424 59051
rect 185264 58989 185424 59023
rect 185264 58961 185299 58989
rect 185327 58961 185361 58989
rect 185389 58961 185424 58989
rect 185264 58944 185424 58961
rect 200624 59175 200784 59192
rect 200624 59147 200659 59175
rect 200687 59147 200721 59175
rect 200749 59147 200784 59175
rect 200624 59113 200784 59147
rect 200624 59085 200659 59113
rect 200687 59085 200721 59113
rect 200749 59085 200784 59113
rect 200624 59051 200784 59085
rect 200624 59023 200659 59051
rect 200687 59023 200721 59051
rect 200749 59023 200784 59051
rect 200624 58989 200784 59023
rect 200624 58961 200659 58989
rect 200687 58961 200721 58989
rect 200749 58961 200784 58989
rect 200624 58944 200784 58961
rect 215984 59175 216144 59192
rect 215984 59147 216019 59175
rect 216047 59147 216081 59175
rect 216109 59147 216144 59175
rect 215984 59113 216144 59147
rect 215984 59085 216019 59113
rect 216047 59085 216081 59113
rect 216109 59085 216144 59113
rect 215984 59051 216144 59085
rect 215984 59023 216019 59051
rect 216047 59023 216081 59051
rect 216109 59023 216144 59051
rect 215984 58989 216144 59023
rect 215984 58961 216019 58989
rect 216047 58961 216081 58989
rect 216109 58961 216144 58989
rect 215984 58944 216144 58961
rect 231344 59175 231504 59192
rect 231344 59147 231379 59175
rect 231407 59147 231441 59175
rect 231469 59147 231504 59175
rect 231344 59113 231504 59147
rect 231344 59085 231379 59113
rect 231407 59085 231441 59113
rect 231469 59085 231504 59113
rect 231344 59051 231504 59085
rect 231344 59023 231379 59051
rect 231407 59023 231441 59051
rect 231469 59023 231504 59051
rect 231344 58989 231504 59023
rect 231344 58961 231379 58989
rect 231407 58961 231441 58989
rect 231469 58961 231504 58989
rect 231344 58944 231504 58961
rect 246704 59175 246864 59192
rect 246704 59147 246739 59175
rect 246767 59147 246801 59175
rect 246829 59147 246864 59175
rect 246704 59113 246864 59147
rect 246704 59085 246739 59113
rect 246767 59085 246801 59113
rect 246829 59085 246864 59113
rect 246704 59051 246864 59085
rect 246704 59023 246739 59051
rect 246767 59023 246801 59051
rect 246829 59023 246864 59051
rect 246704 58989 246864 59023
rect 246704 58961 246739 58989
rect 246767 58961 246801 58989
rect 246829 58961 246864 58989
rect 246704 58944 246864 58961
rect 262064 59175 262224 59192
rect 262064 59147 262099 59175
rect 262127 59147 262161 59175
rect 262189 59147 262224 59175
rect 262064 59113 262224 59147
rect 262064 59085 262099 59113
rect 262127 59085 262161 59113
rect 262189 59085 262224 59113
rect 262064 59051 262224 59085
rect 262064 59023 262099 59051
rect 262127 59023 262161 59051
rect 262189 59023 262224 59051
rect 262064 58989 262224 59023
rect 262064 58961 262099 58989
rect 262127 58961 262161 58989
rect 262189 58961 262224 58989
rect 262064 58944 262224 58961
rect 162224 56175 162384 56192
rect 162224 56147 162259 56175
rect 162287 56147 162321 56175
rect 162349 56147 162384 56175
rect 162224 56113 162384 56147
rect 162224 56085 162259 56113
rect 162287 56085 162321 56113
rect 162349 56085 162384 56113
rect 162224 56051 162384 56085
rect 162224 56023 162259 56051
rect 162287 56023 162321 56051
rect 162349 56023 162384 56051
rect 162224 55989 162384 56023
rect 162224 55961 162259 55989
rect 162287 55961 162321 55989
rect 162349 55961 162384 55989
rect 162224 55944 162384 55961
rect 177584 56175 177744 56192
rect 177584 56147 177619 56175
rect 177647 56147 177681 56175
rect 177709 56147 177744 56175
rect 177584 56113 177744 56147
rect 177584 56085 177619 56113
rect 177647 56085 177681 56113
rect 177709 56085 177744 56113
rect 177584 56051 177744 56085
rect 177584 56023 177619 56051
rect 177647 56023 177681 56051
rect 177709 56023 177744 56051
rect 177584 55989 177744 56023
rect 177584 55961 177619 55989
rect 177647 55961 177681 55989
rect 177709 55961 177744 55989
rect 177584 55944 177744 55961
rect 192944 56175 193104 56192
rect 192944 56147 192979 56175
rect 193007 56147 193041 56175
rect 193069 56147 193104 56175
rect 192944 56113 193104 56147
rect 192944 56085 192979 56113
rect 193007 56085 193041 56113
rect 193069 56085 193104 56113
rect 192944 56051 193104 56085
rect 192944 56023 192979 56051
rect 193007 56023 193041 56051
rect 193069 56023 193104 56051
rect 192944 55989 193104 56023
rect 192944 55961 192979 55989
rect 193007 55961 193041 55989
rect 193069 55961 193104 55989
rect 192944 55944 193104 55961
rect 208304 56175 208464 56192
rect 208304 56147 208339 56175
rect 208367 56147 208401 56175
rect 208429 56147 208464 56175
rect 208304 56113 208464 56147
rect 208304 56085 208339 56113
rect 208367 56085 208401 56113
rect 208429 56085 208464 56113
rect 208304 56051 208464 56085
rect 208304 56023 208339 56051
rect 208367 56023 208401 56051
rect 208429 56023 208464 56051
rect 208304 55989 208464 56023
rect 208304 55961 208339 55989
rect 208367 55961 208401 55989
rect 208429 55961 208464 55989
rect 208304 55944 208464 55961
rect 223664 56175 223824 56192
rect 223664 56147 223699 56175
rect 223727 56147 223761 56175
rect 223789 56147 223824 56175
rect 223664 56113 223824 56147
rect 223664 56085 223699 56113
rect 223727 56085 223761 56113
rect 223789 56085 223824 56113
rect 223664 56051 223824 56085
rect 223664 56023 223699 56051
rect 223727 56023 223761 56051
rect 223789 56023 223824 56051
rect 223664 55989 223824 56023
rect 223664 55961 223699 55989
rect 223727 55961 223761 55989
rect 223789 55961 223824 55989
rect 223664 55944 223824 55961
rect 239024 56175 239184 56192
rect 239024 56147 239059 56175
rect 239087 56147 239121 56175
rect 239149 56147 239184 56175
rect 239024 56113 239184 56147
rect 239024 56085 239059 56113
rect 239087 56085 239121 56113
rect 239149 56085 239184 56113
rect 239024 56051 239184 56085
rect 239024 56023 239059 56051
rect 239087 56023 239121 56051
rect 239149 56023 239184 56051
rect 239024 55989 239184 56023
rect 239024 55961 239059 55989
rect 239087 55961 239121 55989
rect 239149 55961 239184 55989
rect 239024 55944 239184 55961
rect 254384 56175 254544 56192
rect 254384 56147 254419 56175
rect 254447 56147 254481 56175
rect 254509 56147 254544 56175
rect 254384 56113 254544 56147
rect 254384 56085 254419 56113
rect 254447 56085 254481 56113
rect 254509 56085 254544 56113
rect 254384 56051 254544 56085
rect 254384 56023 254419 56051
rect 254447 56023 254481 56051
rect 254509 56023 254544 56051
rect 254384 55989 254544 56023
rect 254384 55961 254419 55989
rect 254447 55961 254481 55989
rect 254509 55961 254544 55989
rect 254384 55944 254544 55961
rect 269744 56175 269904 56192
rect 269744 56147 269779 56175
rect 269807 56147 269841 56175
rect 269869 56147 269904 56175
rect 269744 56113 269904 56147
rect 269744 56085 269779 56113
rect 269807 56085 269841 56113
rect 269869 56085 269904 56113
rect 269744 56051 269904 56085
rect 269744 56023 269779 56051
rect 269807 56023 269841 56051
rect 269869 56023 269904 56051
rect 269744 55989 269904 56023
rect 269744 55961 269779 55989
rect 269807 55961 269841 55989
rect 269869 55961 269904 55989
rect 269744 55944 269904 55961
rect 158169 50147 158217 50175
rect 158245 50147 158279 50175
rect 158307 50147 158341 50175
rect 158369 50147 158403 50175
rect 158431 50147 158479 50175
rect 158169 50113 158479 50147
rect 158169 50085 158217 50113
rect 158245 50085 158279 50113
rect 158307 50085 158341 50113
rect 158369 50085 158403 50113
rect 158431 50085 158479 50113
rect 158169 50051 158479 50085
rect 158169 50023 158217 50051
rect 158245 50023 158279 50051
rect 158307 50023 158341 50051
rect 158369 50023 158403 50051
rect 158431 50023 158479 50051
rect 158169 49989 158479 50023
rect 158169 49961 158217 49989
rect 158245 49961 158279 49989
rect 158307 49961 158341 49989
rect 158369 49961 158403 49989
rect 158431 49961 158479 49989
rect 158169 41175 158479 49961
rect 169904 50175 170064 50192
rect 169904 50147 169939 50175
rect 169967 50147 170001 50175
rect 170029 50147 170064 50175
rect 169904 50113 170064 50147
rect 169904 50085 169939 50113
rect 169967 50085 170001 50113
rect 170029 50085 170064 50113
rect 169904 50051 170064 50085
rect 169904 50023 169939 50051
rect 169967 50023 170001 50051
rect 170029 50023 170064 50051
rect 169904 49989 170064 50023
rect 169904 49961 169939 49989
rect 169967 49961 170001 49989
rect 170029 49961 170064 49989
rect 169904 49944 170064 49961
rect 185264 50175 185424 50192
rect 185264 50147 185299 50175
rect 185327 50147 185361 50175
rect 185389 50147 185424 50175
rect 185264 50113 185424 50147
rect 185264 50085 185299 50113
rect 185327 50085 185361 50113
rect 185389 50085 185424 50113
rect 185264 50051 185424 50085
rect 185264 50023 185299 50051
rect 185327 50023 185361 50051
rect 185389 50023 185424 50051
rect 185264 49989 185424 50023
rect 185264 49961 185299 49989
rect 185327 49961 185361 49989
rect 185389 49961 185424 49989
rect 185264 49944 185424 49961
rect 200624 50175 200784 50192
rect 200624 50147 200659 50175
rect 200687 50147 200721 50175
rect 200749 50147 200784 50175
rect 200624 50113 200784 50147
rect 200624 50085 200659 50113
rect 200687 50085 200721 50113
rect 200749 50085 200784 50113
rect 200624 50051 200784 50085
rect 200624 50023 200659 50051
rect 200687 50023 200721 50051
rect 200749 50023 200784 50051
rect 200624 49989 200784 50023
rect 200624 49961 200659 49989
rect 200687 49961 200721 49989
rect 200749 49961 200784 49989
rect 200624 49944 200784 49961
rect 215984 50175 216144 50192
rect 215984 50147 216019 50175
rect 216047 50147 216081 50175
rect 216109 50147 216144 50175
rect 215984 50113 216144 50147
rect 215984 50085 216019 50113
rect 216047 50085 216081 50113
rect 216109 50085 216144 50113
rect 215984 50051 216144 50085
rect 215984 50023 216019 50051
rect 216047 50023 216081 50051
rect 216109 50023 216144 50051
rect 215984 49989 216144 50023
rect 215984 49961 216019 49989
rect 216047 49961 216081 49989
rect 216109 49961 216144 49989
rect 215984 49944 216144 49961
rect 231344 50175 231504 50192
rect 231344 50147 231379 50175
rect 231407 50147 231441 50175
rect 231469 50147 231504 50175
rect 231344 50113 231504 50147
rect 231344 50085 231379 50113
rect 231407 50085 231441 50113
rect 231469 50085 231504 50113
rect 231344 50051 231504 50085
rect 231344 50023 231379 50051
rect 231407 50023 231441 50051
rect 231469 50023 231504 50051
rect 231344 49989 231504 50023
rect 231344 49961 231379 49989
rect 231407 49961 231441 49989
rect 231469 49961 231504 49989
rect 231344 49944 231504 49961
rect 246704 50175 246864 50192
rect 246704 50147 246739 50175
rect 246767 50147 246801 50175
rect 246829 50147 246864 50175
rect 246704 50113 246864 50147
rect 246704 50085 246739 50113
rect 246767 50085 246801 50113
rect 246829 50085 246864 50113
rect 246704 50051 246864 50085
rect 246704 50023 246739 50051
rect 246767 50023 246801 50051
rect 246829 50023 246864 50051
rect 246704 49989 246864 50023
rect 246704 49961 246739 49989
rect 246767 49961 246801 49989
rect 246829 49961 246864 49989
rect 246704 49944 246864 49961
rect 262064 50175 262224 50192
rect 262064 50147 262099 50175
rect 262127 50147 262161 50175
rect 262189 50147 262224 50175
rect 262064 50113 262224 50147
rect 262064 50085 262099 50113
rect 262127 50085 262161 50113
rect 262189 50085 262224 50113
rect 262064 50051 262224 50085
rect 262064 50023 262099 50051
rect 262127 50023 262161 50051
rect 262189 50023 262224 50051
rect 262064 49989 262224 50023
rect 262064 49961 262099 49989
rect 262127 49961 262161 49989
rect 262189 49961 262224 49989
rect 262064 49944 262224 49961
rect 162224 47175 162384 47192
rect 162224 47147 162259 47175
rect 162287 47147 162321 47175
rect 162349 47147 162384 47175
rect 162224 47113 162384 47147
rect 162224 47085 162259 47113
rect 162287 47085 162321 47113
rect 162349 47085 162384 47113
rect 162224 47051 162384 47085
rect 162224 47023 162259 47051
rect 162287 47023 162321 47051
rect 162349 47023 162384 47051
rect 162224 46989 162384 47023
rect 162224 46961 162259 46989
rect 162287 46961 162321 46989
rect 162349 46961 162384 46989
rect 162224 46944 162384 46961
rect 177584 47175 177744 47192
rect 177584 47147 177619 47175
rect 177647 47147 177681 47175
rect 177709 47147 177744 47175
rect 177584 47113 177744 47147
rect 177584 47085 177619 47113
rect 177647 47085 177681 47113
rect 177709 47085 177744 47113
rect 177584 47051 177744 47085
rect 177584 47023 177619 47051
rect 177647 47023 177681 47051
rect 177709 47023 177744 47051
rect 177584 46989 177744 47023
rect 177584 46961 177619 46989
rect 177647 46961 177681 46989
rect 177709 46961 177744 46989
rect 177584 46944 177744 46961
rect 192944 47175 193104 47192
rect 192944 47147 192979 47175
rect 193007 47147 193041 47175
rect 193069 47147 193104 47175
rect 192944 47113 193104 47147
rect 192944 47085 192979 47113
rect 193007 47085 193041 47113
rect 193069 47085 193104 47113
rect 192944 47051 193104 47085
rect 192944 47023 192979 47051
rect 193007 47023 193041 47051
rect 193069 47023 193104 47051
rect 192944 46989 193104 47023
rect 192944 46961 192979 46989
rect 193007 46961 193041 46989
rect 193069 46961 193104 46989
rect 192944 46944 193104 46961
rect 208304 47175 208464 47192
rect 208304 47147 208339 47175
rect 208367 47147 208401 47175
rect 208429 47147 208464 47175
rect 208304 47113 208464 47147
rect 208304 47085 208339 47113
rect 208367 47085 208401 47113
rect 208429 47085 208464 47113
rect 208304 47051 208464 47085
rect 208304 47023 208339 47051
rect 208367 47023 208401 47051
rect 208429 47023 208464 47051
rect 208304 46989 208464 47023
rect 208304 46961 208339 46989
rect 208367 46961 208401 46989
rect 208429 46961 208464 46989
rect 208304 46944 208464 46961
rect 223664 47175 223824 47192
rect 223664 47147 223699 47175
rect 223727 47147 223761 47175
rect 223789 47147 223824 47175
rect 223664 47113 223824 47147
rect 223664 47085 223699 47113
rect 223727 47085 223761 47113
rect 223789 47085 223824 47113
rect 223664 47051 223824 47085
rect 223664 47023 223699 47051
rect 223727 47023 223761 47051
rect 223789 47023 223824 47051
rect 223664 46989 223824 47023
rect 223664 46961 223699 46989
rect 223727 46961 223761 46989
rect 223789 46961 223824 46989
rect 223664 46944 223824 46961
rect 239024 47175 239184 47192
rect 239024 47147 239059 47175
rect 239087 47147 239121 47175
rect 239149 47147 239184 47175
rect 239024 47113 239184 47147
rect 239024 47085 239059 47113
rect 239087 47085 239121 47113
rect 239149 47085 239184 47113
rect 239024 47051 239184 47085
rect 239024 47023 239059 47051
rect 239087 47023 239121 47051
rect 239149 47023 239184 47051
rect 239024 46989 239184 47023
rect 239024 46961 239059 46989
rect 239087 46961 239121 46989
rect 239149 46961 239184 46989
rect 239024 46944 239184 46961
rect 254384 47175 254544 47192
rect 254384 47147 254419 47175
rect 254447 47147 254481 47175
rect 254509 47147 254544 47175
rect 254384 47113 254544 47147
rect 254384 47085 254419 47113
rect 254447 47085 254481 47113
rect 254509 47085 254544 47113
rect 254384 47051 254544 47085
rect 254384 47023 254419 47051
rect 254447 47023 254481 47051
rect 254509 47023 254544 47051
rect 254384 46989 254544 47023
rect 254384 46961 254419 46989
rect 254447 46961 254481 46989
rect 254509 46961 254544 46989
rect 254384 46944 254544 46961
rect 269744 47175 269904 47192
rect 269744 47147 269779 47175
rect 269807 47147 269841 47175
rect 269869 47147 269904 47175
rect 269744 47113 269904 47147
rect 269744 47085 269779 47113
rect 269807 47085 269841 47113
rect 269869 47085 269904 47113
rect 269744 47051 269904 47085
rect 269744 47023 269779 47051
rect 269807 47023 269841 47051
rect 269869 47023 269904 47051
rect 269744 46989 269904 47023
rect 269744 46961 269779 46989
rect 269807 46961 269841 46989
rect 269869 46961 269904 46989
rect 269744 46944 269904 46961
rect 158169 41147 158217 41175
rect 158245 41147 158279 41175
rect 158307 41147 158341 41175
rect 158369 41147 158403 41175
rect 158431 41147 158479 41175
rect 158169 41113 158479 41147
rect 158169 41085 158217 41113
rect 158245 41085 158279 41113
rect 158307 41085 158341 41113
rect 158369 41085 158403 41113
rect 158431 41085 158479 41113
rect 158169 41051 158479 41085
rect 158169 41023 158217 41051
rect 158245 41023 158279 41051
rect 158307 41023 158341 41051
rect 158369 41023 158403 41051
rect 158431 41023 158479 41051
rect 158169 40989 158479 41023
rect 158169 40961 158217 40989
rect 158245 40961 158279 40989
rect 158307 40961 158341 40989
rect 158369 40961 158403 40989
rect 158431 40961 158479 40989
rect 158169 32175 158479 40961
rect 169904 41175 170064 41192
rect 169904 41147 169939 41175
rect 169967 41147 170001 41175
rect 170029 41147 170064 41175
rect 169904 41113 170064 41147
rect 169904 41085 169939 41113
rect 169967 41085 170001 41113
rect 170029 41085 170064 41113
rect 169904 41051 170064 41085
rect 169904 41023 169939 41051
rect 169967 41023 170001 41051
rect 170029 41023 170064 41051
rect 169904 40989 170064 41023
rect 169904 40961 169939 40989
rect 169967 40961 170001 40989
rect 170029 40961 170064 40989
rect 169904 40944 170064 40961
rect 185264 41175 185424 41192
rect 185264 41147 185299 41175
rect 185327 41147 185361 41175
rect 185389 41147 185424 41175
rect 185264 41113 185424 41147
rect 185264 41085 185299 41113
rect 185327 41085 185361 41113
rect 185389 41085 185424 41113
rect 185264 41051 185424 41085
rect 185264 41023 185299 41051
rect 185327 41023 185361 41051
rect 185389 41023 185424 41051
rect 185264 40989 185424 41023
rect 185264 40961 185299 40989
rect 185327 40961 185361 40989
rect 185389 40961 185424 40989
rect 185264 40944 185424 40961
rect 200624 41175 200784 41192
rect 200624 41147 200659 41175
rect 200687 41147 200721 41175
rect 200749 41147 200784 41175
rect 200624 41113 200784 41147
rect 200624 41085 200659 41113
rect 200687 41085 200721 41113
rect 200749 41085 200784 41113
rect 200624 41051 200784 41085
rect 200624 41023 200659 41051
rect 200687 41023 200721 41051
rect 200749 41023 200784 41051
rect 200624 40989 200784 41023
rect 200624 40961 200659 40989
rect 200687 40961 200721 40989
rect 200749 40961 200784 40989
rect 200624 40944 200784 40961
rect 215984 41175 216144 41192
rect 215984 41147 216019 41175
rect 216047 41147 216081 41175
rect 216109 41147 216144 41175
rect 215984 41113 216144 41147
rect 215984 41085 216019 41113
rect 216047 41085 216081 41113
rect 216109 41085 216144 41113
rect 215984 41051 216144 41085
rect 215984 41023 216019 41051
rect 216047 41023 216081 41051
rect 216109 41023 216144 41051
rect 215984 40989 216144 41023
rect 215984 40961 216019 40989
rect 216047 40961 216081 40989
rect 216109 40961 216144 40989
rect 215984 40944 216144 40961
rect 231344 41175 231504 41192
rect 231344 41147 231379 41175
rect 231407 41147 231441 41175
rect 231469 41147 231504 41175
rect 231344 41113 231504 41147
rect 231344 41085 231379 41113
rect 231407 41085 231441 41113
rect 231469 41085 231504 41113
rect 231344 41051 231504 41085
rect 231344 41023 231379 41051
rect 231407 41023 231441 41051
rect 231469 41023 231504 41051
rect 231344 40989 231504 41023
rect 231344 40961 231379 40989
rect 231407 40961 231441 40989
rect 231469 40961 231504 40989
rect 231344 40944 231504 40961
rect 246704 41175 246864 41192
rect 246704 41147 246739 41175
rect 246767 41147 246801 41175
rect 246829 41147 246864 41175
rect 246704 41113 246864 41147
rect 246704 41085 246739 41113
rect 246767 41085 246801 41113
rect 246829 41085 246864 41113
rect 246704 41051 246864 41085
rect 246704 41023 246739 41051
rect 246767 41023 246801 41051
rect 246829 41023 246864 41051
rect 246704 40989 246864 41023
rect 246704 40961 246739 40989
rect 246767 40961 246801 40989
rect 246829 40961 246864 40989
rect 246704 40944 246864 40961
rect 262064 41175 262224 41192
rect 262064 41147 262099 41175
rect 262127 41147 262161 41175
rect 262189 41147 262224 41175
rect 262064 41113 262224 41147
rect 262064 41085 262099 41113
rect 262127 41085 262161 41113
rect 262189 41085 262224 41113
rect 262064 41051 262224 41085
rect 262064 41023 262099 41051
rect 262127 41023 262161 41051
rect 262189 41023 262224 41051
rect 262064 40989 262224 41023
rect 262064 40961 262099 40989
rect 262127 40961 262161 40989
rect 262189 40961 262224 40989
rect 262064 40944 262224 40961
rect 162224 38175 162384 38192
rect 162224 38147 162259 38175
rect 162287 38147 162321 38175
rect 162349 38147 162384 38175
rect 162224 38113 162384 38147
rect 162224 38085 162259 38113
rect 162287 38085 162321 38113
rect 162349 38085 162384 38113
rect 162224 38051 162384 38085
rect 162224 38023 162259 38051
rect 162287 38023 162321 38051
rect 162349 38023 162384 38051
rect 162224 37989 162384 38023
rect 162224 37961 162259 37989
rect 162287 37961 162321 37989
rect 162349 37961 162384 37989
rect 162224 37944 162384 37961
rect 177584 38175 177744 38192
rect 177584 38147 177619 38175
rect 177647 38147 177681 38175
rect 177709 38147 177744 38175
rect 177584 38113 177744 38147
rect 177584 38085 177619 38113
rect 177647 38085 177681 38113
rect 177709 38085 177744 38113
rect 177584 38051 177744 38085
rect 177584 38023 177619 38051
rect 177647 38023 177681 38051
rect 177709 38023 177744 38051
rect 177584 37989 177744 38023
rect 177584 37961 177619 37989
rect 177647 37961 177681 37989
rect 177709 37961 177744 37989
rect 177584 37944 177744 37961
rect 192944 38175 193104 38192
rect 192944 38147 192979 38175
rect 193007 38147 193041 38175
rect 193069 38147 193104 38175
rect 192944 38113 193104 38147
rect 192944 38085 192979 38113
rect 193007 38085 193041 38113
rect 193069 38085 193104 38113
rect 192944 38051 193104 38085
rect 192944 38023 192979 38051
rect 193007 38023 193041 38051
rect 193069 38023 193104 38051
rect 192944 37989 193104 38023
rect 192944 37961 192979 37989
rect 193007 37961 193041 37989
rect 193069 37961 193104 37989
rect 192944 37944 193104 37961
rect 208304 38175 208464 38192
rect 208304 38147 208339 38175
rect 208367 38147 208401 38175
rect 208429 38147 208464 38175
rect 208304 38113 208464 38147
rect 208304 38085 208339 38113
rect 208367 38085 208401 38113
rect 208429 38085 208464 38113
rect 208304 38051 208464 38085
rect 208304 38023 208339 38051
rect 208367 38023 208401 38051
rect 208429 38023 208464 38051
rect 208304 37989 208464 38023
rect 208304 37961 208339 37989
rect 208367 37961 208401 37989
rect 208429 37961 208464 37989
rect 208304 37944 208464 37961
rect 223664 38175 223824 38192
rect 223664 38147 223699 38175
rect 223727 38147 223761 38175
rect 223789 38147 223824 38175
rect 223664 38113 223824 38147
rect 223664 38085 223699 38113
rect 223727 38085 223761 38113
rect 223789 38085 223824 38113
rect 223664 38051 223824 38085
rect 223664 38023 223699 38051
rect 223727 38023 223761 38051
rect 223789 38023 223824 38051
rect 223664 37989 223824 38023
rect 223664 37961 223699 37989
rect 223727 37961 223761 37989
rect 223789 37961 223824 37989
rect 223664 37944 223824 37961
rect 239024 38175 239184 38192
rect 239024 38147 239059 38175
rect 239087 38147 239121 38175
rect 239149 38147 239184 38175
rect 239024 38113 239184 38147
rect 239024 38085 239059 38113
rect 239087 38085 239121 38113
rect 239149 38085 239184 38113
rect 239024 38051 239184 38085
rect 239024 38023 239059 38051
rect 239087 38023 239121 38051
rect 239149 38023 239184 38051
rect 239024 37989 239184 38023
rect 239024 37961 239059 37989
rect 239087 37961 239121 37989
rect 239149 37961 239184 37989
rect 239024 37944 239184 37961
rect 254384 38175 254544 38192
rect 254384 38147 254419 38175
rect 254447 38147 254481 38175
rect 254509 38147 254544 38175
rect 254384 38113 254544 38147
rect 254384 38085 254419 38113
rect 254447 38085 254481 38113
rect 254509 38085 254544 38113
rect 254384 38051 254544 38085
rect 254384 38023 254419 38051
rect 254447 38023 254481 38051
rect 254509 38023 254544 38051
rect 254384 37989 254544 38023
rect 254384 37961 254419 37989
rect 254447 37961 254481 37989
rect 254509 37961 254544 37989
rect 254384 37944 254544 37961
rect 269744 38175 269904 38192
rect 269744 38147 269779 38175
rect 269807 38147 269841 38175
rect 269869 38147 269904 38175
rect 269744 38113 269904 38147
rect 269744 38085 269779 38113
rect 269807 38085 269841 38113
rect 269869 38085 269904 38113
rect 269744 38051 269904 38085
rect 269744 38023 269779 38051
rect 269807 38023 269841 38051
rect 269869 38023 269904 38051
rect 269744 37989 269904 38023
rect 269744 37961 269779 37989
rect 269807 37961 269841 37989
rect 269869 37961 269904 37989
rect 269744 37944 269904 37961
rect 158169 32147 158217 32175
rect 158245 32147 158279 32175
rect 158307 32147 158341 32175
rect 158369 32147 158403 32175
rect 158431 32147 158479 32175
rect 158169 32113 158479 32147
rect 158169 32085 158217 32113
rect 158245 32085 158279 32113
rect 158307 32085 158341 32113
rect 158369 32085 158403 32113
rect 158431 32085 158479 32113
rect 158169 32051 158479 32085
rect 158169 32023 158217 32051
rect 158245 32023 158279 32051
rect 158307 32023 158341 32051
rect 158369 32023 158403 32051
rect 158431 32023 158479 32051
rect 158169 31989 158479 32023
rect 158169 31961 158217 31989
rect 158245 31961 158279 31989
rect 158307 31961 158341 31989
rect 158369 31961 158403 31989
rect 158431 31961 158479 31989
rect 158169 23175 158479 31961
rect 169904 32175 170064 32192
rect 169904 32147 169939 32175
rect 169967 32147 170001 32175
rect 170029 32147 170064 32175
rect 169904 32113 170064 32147
rect 169904 32085 169939 32113
rect 169967 32085 170001 32113
rect 170029 32085 170064 32113
rect 169904 32051 170064 32085
rect 169904 32023 169939 32051
rect 169967 32023 170001 32051
rect 170029 32023 170064 32051
rect 169904 31989 170064 32023
rect 169904 31961 169939 31989
rect 169967 31961 170001 31989
rect 170029 31961 170064 31989
rect 169904 31944 170064 31961
rect 185264 32175 185424 32192
rect 185264 32147 185299 32175
rect 185327 32147 185361 32175
rect 185389 32147 185424 32175
rect 185264 32113 185424 32147
rect 185264 32085 185299 32113
rect 185327 32085 185361 32113
rect 185389 32085 185424 32113
rect 185264 32051 185424 32085
rect 185264 32023 185299 32051
rect 185327 32023 185361 32051
rect 185389 32023 185424 32051
rect 185264 31989 185424 32023
rect 185264 31961 185299 31989
rect 185327 31961 185361 31989
rect 185389 31961 185424 31989
rect 185264 31944 185424 31961
rect 200624 32175 200784 32192
rect 200624 32147 200659 32175
rect 200687 32147 200721 32175
rect 200749 32147 200784 32175
rect 200624 32113 200784 32147
rect 200624 32085 200659 32113
rect 200687 32085 200721 32113
rect 200749 32085 200784 32113
rect 200624 32051 200784 32085
rect 200624 32023 200659 32051
rect 200687 32023 200721 32051
rect 200749 32023 200784 32051
rect 200624 31989 200784 32023
rect 200624 31961 200659 31989
rect 200687 31961 200721 31989
rect 200749 31961 200784 31989
rect 200624 31944 200784 31961
rect 215984 32175 216144 32192
rect 215984 32147 216019 32175
rect 216047 32147 216081 32175
rect 216109 32147 216144 32175
rect 215984 32113 216144 32147
rect 215984 32085 216019 32113
rect 216047 32085 216081 32113
rect 216109 32085 216144 32113
rect 215984 32051 216144 32085
rect 215984 32023 216019 32051
rect 216047 32023 216081 32051
rect 216109 32023 216144 32051
rect 215984 31989 216144 32023
rect 215984 31961 216019 31989
rect 216047 31961 216081 31989
rect 216109 31961 216144 31989
rect 215984 31944 216144 31961
rect 231344 32175 231504 32192
rect 231344 32147 231379 32175
rect 231407 32147 231441 32175
rect 231469 32147 231504 32175
rect 231344 32113 231504 32147
rect 231344 32085 231379 32113
rect 231407 32085 231441 32113
rect 231469 32085 231504 32113
rect 231344 32051 231504 32085
rect 231344 32023 231379 32051
rect 231407 32023 231441 32051
rect 231469 32023 231504 32051
rect 231344 31989 231504 32023
rect 231344 31961 231379 31989
rect 231407 31961 231441 31989
rect 231469 31961 231504 31989
rect 231344 31944 231504 31961
rect 246704 32175 246864 32192
rect 246704 32147 246739 32175
rect 246767 32147 246801 32175
rect 246829 32147 246864 32175
rect 246704 32113 246864 32147
rect 246704 32085 246739 32113
rect 246767 32085 246801 32113
rect 246829 32085 246864 32113
rect 246704 32051 246864 32085
rect 246704 32023 246739 32051
rect 246767 32023 246801 32051
rect 246829 32023 246864 32051
rect 246704 31989 246864 32023
rect 246704 31961 246739 31989
rect 246767 31961 246801 31989
rect 246829 31961 246864 31989
rect 246704 31944 246864 31961
rect 262064 32175 262224 32192
rect 262064 32147 262099 32175
rect 262127 32147 262161 32175
rect 262189 32147 262224 32175
rect 262064 32113 262224 32147
rect 262064 32085 262099 32113
rect 262127 32085 262161 32113
rect 262189 32085 262224 32113
rect 262064 32051 262224 32085
rect 262064 32023 262099 32051
rect 262127 32023 262161 32051
rect 262189 32023 262224 32051
rect 262064 31989 262224 32023
rect 262064 31961 262099 31989
rect 262127 31961 262161 31989
rect 262189 31961 262224 31989
rect 262064 31944 262224 31961
rect 162224 29175 162384 29192
rect 162224 29147 162259 29175
rect 162287 29147 162321 29175
rect 162349 29147 162384 29175
rect 162224 29113 162384 29147
rect 162224 29085 162259 29113
rect 162287 29085 162321 29113
rect 162349 29085 162384 29113
rect 162224 29051 162384 29085
rect 162224 29023 162259 29051
rect 162287 29023 162321 29051
rect 162349 29023 162384 29051
rect 162224 28989 162384 29023
rect 162224 28961 162259 28989
rect 162287 28961 162321 28989
rect 162349 28961 162384 28989
rect 162224 28944 162384 28961
rect 177584 29175 177744 29192
rect 177584 29147 177619 29175
rect 177647 29147 177681 29175
rect 177709 29147 177744 29175
rect 177584 29113 177744 29147
rect 177584 29085 177619 29113
rect 177647 29085 177681 29113
rect 177709 29085 177744 29113
rect 177584 29051 177744 29085
rect 177584 29023 177619 29051
rect 177647 29023 177681 29051
rect 177709 29023 177744 29051
rect 177584 28989 177744 29023
rect 177584 28961 177619 28989
rect 177647 28961 177681 28989
rect 177709 28961 177744 28989
rect 177584 28944 177744 28961
rect 192944 29175 193104 29192
rect 192944 29147 192979 29175
rect 193007 29147 193041 29175
rect 193069 29147 193104 29175
rect 192944 29113 193104 29147
rect 192944 29085 192979 29113
rect 193007 29085 193041 29113
rect 193069 29085 193104 29113
rect 192944 29051 193104 29085
rect 192944 29023 192979 29051
rect 193007 29023 193041 29051
rect 193069 29023 193104 29051
rect 192944 28989 193104 29023
rect 192944 28961 192979 28989
rect 193007 28961 193041 28989
rect 193069 28961 193104 28989
rect 192944 28944 193104 28961
rect 208304 29175 208464 29192
rect 208304 29147 208339 29175
rect 208367 29147 208401 29175
rect 208429 29147 208464 29175
rect 208304 29113 208464 29147
rect 208304 29085 208339 29113
rect 208367 29085 208401 29113
rect 208429 29085 208464 29113
rect 208304 29051 208464 29085
rect 208304 29023 208339 29051
rect 208367 29023 208401 29051
rect 208429 29023 208464 29051
rect 208304 28989 208464 29023
rect 208304 28961 208339 28989
rect 208367 28961 208401 28989
rect 208429 28961 208464 28989
rect 208304 28944 208464 28961
rect 223664 29175 223824 29192
rect 223664 29147 223699 29175
rect 223727 29147 223761 29175
rect 223789 29147 223824 29175
rect 223664 29113 223824 29147
rect 223664 29085 223699 29113
rect 223727 29085 223761 29113
rect 223789 29085 223824 29113
rect 223664 29051 223824 29085
rect 223664 29023 223699 29051
rect 223727 29023 223761 29051
rect 223789 29023 223824 29051
rect 223664 28989 223824 29023
rect 223664 28961 223699 28989
rect 223727 28961 223761 28989
rect 223789 28961 223824 28989
rect 223664 28944 223824 28961
rect 239024 29175 239184 29192
rect 239024 29147 239059 29175
rect 239087 29147 239121 29175
rect 239149 29147 239184 29175
rect 239024 29113 239184 29147
rect 239024 29085 239059 29113
rect 239087 29085 239121 29113
rect 239149 29085 239184 29113
rect 239024 29051 239184 29085
rect 239024 29023 239059 29051
rect 239087 29023 239121 29051
rect 239149 29023 239184 29051
rect 239024 28989 239184 29023
rect 239024 28961 239059 28989
rect 239087 28961 239121 28989
rect 239149 28961 239184 28989
rect 239024 28944 239184 28961
rect 254384 29175 254544 29192
rect 254384 29147 254419 29175
rect 254447 29147 254481 29175
rect 254509 29147 254544 29175
rect 254384 29113 254544 29147
rect 254384 29085 254419 29113
rect 254447 29085 254481 29113
rect 254509 29085 254544 29113
rect 254384 29051 254544 29085
rect 254384 29023 254419 29051
rect 254447 29023 254481 29051
rect 254509 29023 254544 29051
rect 254384 28989 254544 29023
rect 254384 28961 254419 28989
rect 254447 28961 254481 28989
rect 254509 28961 254544 28989
rect 254384 28944 254544 28961
rect 269744 29175 269904 29192
rect 269744 29147 269779 29175
rect 269807 29147 269841 29175
rect 269869 29147 269904 29175
rect 269744 29113 269904 29147
rect 269744 29085 269779 29113
rect 269807 29085 269841 29113
rect 269869 29085 269904 29113
rect 269744 29051 269904 29085
rect 269744 29023 269779 29051
rect 269807 29023 269841 29051
rect 269869 29023 269904 29051
rect 269744 28989 269904 29023
rect 269744 28961 269779 28989
rect 269807 28961 269841 28989
rect 269869 28961 269904 28989
rect 269744 28944 269904 28961
rect 158169 23147 158217 23175
rect 158245 23147 158279 23175
rect 158307 23147 158341 23175
rect 158369 23147 158403 23175
rect 158431 23147 158479 23175
rect 158169 23113 158479 23147
rect 158169 23085 158217 23113
rect 158245 23085 158279 23113
rect 158307 23085 158341 23113
rect 158369 23085 158403 23113
rect 158431 23085 158479 23113
rect 158169 23051 158479 23085
rect 158169 23023 158217 23051
rect 158245 23023 158279 23051
rect 158307 23023 158341 23051
rect 158369 23023 158403 23051
rect 158431 23023 158479 23051
rect 158169 22989 158479 23023
rect 158169 22961 158217 22989
rect 158245 22961 158279 22989
rect 158307 22961 158341 22989
rect 158369 22961 158403 22989
rect 158431 22961 158479 22989
rect 158169 14175 158479 22961
rect 169904 23175 170064 23192
rect 169904 23147 169939 23175
rect 169967 23147 170001 23175
rect 170029 23147 170064 23175
rect 169904 23113 170064 23147
rect 169904 23085 169939 23113
rect 169967 23085 170001 23113
rect 170029 23085 170064 23113
rect 169904 23051 170064 23085
rect 169904 23023 169939 23051
rect 169967 23023 170001 23051
rect 170029 23023 170064 23051
rect 169904 22989 170064 23023
rect 169904 22961 169939 22989
rect 169967 22961 170001 22989
rect 170029 22961 170064 22989
rect 169904 22944 170064 22961
rect 185264 23175 185424 23192
rect 185264 23147 185299 23175
rect 185327 23147 185361 23175
rect 185389 23147 185424 23175
rect 185264 23113 185424 23147
rect 185264 23085 185299 23113
rect 185327 23085 185361 23113
rect 185389 23085 185424 23113
rect 185264 23051 185424 23085
rect 185264 23023 185299 23051
rect 185327 23023 185361 23051
rect 185389 23023 185424 23051
rect 185264 22989 185424 23023
rect 185264 22961 185299 22989
rect 185327 22961 185361 22989
rect 185389 22961 185424 22989
rect 185264 22944 185424 22961
rect 200624 23175 200784 23192
rect 200624 23147 200659 23175
rect 200687 23147 200721 23175
rect 200749 23147 200784 23175
rect 200624 23113 200784 23147
rect 200624 23085 200659 23113
rect 200687 23085 200721 23113
rect 200749 23085 200784 23113
rect 200624 23051 200784 23085
rect 200624 23023 200659 23051
rect 200687 23023 200721 23051
rect 200749 23023 200784 23051
rect 200624 22989 200784 23023
rect 200624 22961 200659 22989
rect 200687 22961 200721 22989
rect 200749 22961 200784 22989
rect 200624 22944 200784 22961
rect 215984 23175 216144 23192
rect 215984 23147 216019 23175
rect 216047 23147 216081 23175
rect 216109 23147 216144 23175
rect 215984 23113 216144 23147
rect 215984 23085 216019 23113
rect 216047 23085 216081 23113
rect 216109 23085 216144 23113
rect 215984 23051 216144 23085
rect 215984 23023 216019 23051
rect 216047 23023 216081 23051
rect 216109 23023 216144 23051
rect 215984 22989 216144 23023
rect 215984 22961 216019 22989
rect 216047 22961 216081 22989
rect 216109 22961 216144 22989
rect 215984 22944 216144 22961
rect 231344 23175 231504 23192
rect 231344 23147 231379 23175
rect 231407 23147 231441 23175
rect 231469 23147 231504 23175
rect 231344 23113 231504 23147
rect 231344 23085 231379 23113
rect 231407 23085 231441 23113
rect 231469 23085 231504 23113
rect 231344 23051 231504 23085
rect 231344 23023 231379 23051
rect 231407 23023 231441 23051
rect 231469 23023 231504 23051
rect 231344 22989 231504 23023
rect 231344 22961 231379 22989
rect 231407 22961 231441 22989
rect 231469 22961 231504 22989
rect 231344 22944 231504 22961
rect 246704 23175 246864 23192
rect 246704 23147 246739 23175
rect 246767 23147 246801 23175
rect 246829 23147 246864 23175
rect 246704 23113 246864 23147
rect 246704 23085 246739 23113
rect 246767 23085 246801 23113
rect 246829 23085 246864 23113
rect 246704 23051 246864 23085
rect 246704 23023 246739 23051
rect 246767 23023 246801 23051
rect 246829 23023 246864 23051
rect 246704 22989 246864 23023
rect 246704 22961 246739 22989
rect 246767 22961 246801 22989
rect 246829 22961 246864 22989
rect 246704 22944 246864 22961
rect 262064 23175 262224 23192
rect 262064 23147 262099 23175
rect 262127 23147 262161 23175
rect 262189 23147 262224 23175
rect 262064 23113 262224 23147
rect 262064 23085 262099 23113
rect 262127 23085 262161 23113
rect 262189 23085 262224 23113
rect 262064 23051 262224 23085
rect 262064 23023 262099 23051
rect 262127 23023 262161 23051
rect 262189 23023 262224 23051
rect 262064 22989 262224 23023
rect 262064 22961 262099 22989
rect 262127 22961 262161 22989
rect 262189 22961 262224 22989
rect 262064 22944 262224 22961
rect 162224 20175 162384 20192
rect 162224 20147 162259 20175
rect 162287 20147 162321 20175
rect 162349 20147 162384 20175
rect 162224 20113 162384 20147
rect 162224 20085 162259 20113
rect 162287 20085 162321 20113
rect 162349 20085 162384 20113
rect 162224 20051 162384 20085
rect 162224 20023 162259 20051
rect 162287 20023 162321 20051
rect 162349 20023 162384 20051
rect 162224 19989 162384 20023
rect 162224 19961 162259 19989
rect 162287 19961 162321 19989
rect 162349 19961 162384 19989
rect 162224 19944 162384 19961
rect 177584 20175 177744 20192
rect 177584 20147 177619 20175
rect 177647 20147 177681 20175
rect 177709 20147 177744 20175
rect 177584 20113 177744 20147
rect 177584 20085 177619 20113
rect 177647 20085 177681 20113
rect 177709 20085 177744 20113
rect 177584 20051 177744 20085
rect 177584 20023 177619 20051
rect 177647 20023 177681 20051
rect 177709 20023 177744 20051
rect 177584 19989 177744 20023
rect 177584 19961 177619 19989
rect 177647 19961 177681 19989
rect 177709 19961 177744 19989
rect 177584 19944 177744 19961
rect 192944 20175 193104 20192
rect 192944 20147 192979 20175
rect 193007 20147 193041 20175
rect 193069 20147 193104 20175
rect 192944 20113 193104 20147
rect 192944 20085 192979 20113
rect 193007 20085 193041 20113
rect 193069 20085 193104 20113
rect 192944 20051 193104 20085
rect 192944 20023 192979 20051
rect 193007 20023 193041 20051
rect 193069 20023 193104 20051
rect 192944 19989 193104 20023
rect 192944 19961 192979 19989
rect 193007 19961 193041 19989
rect 193069 19961 193104 19989
rect 192944 19944 193104 19961
rect 208304 20175 208464 20192
rect 208304 20147 208339 20175
rect 208367 20147 208401 20175
rect 208429 20147 208464 20175
rect 208304 20113 208464 20147
rect 208304 20085 208339 20113
rect 208367 20085 208401 20113
rect 208429 20085 208464 20113
rect 208304 20051 208464 20085
rect 208304 20023 208339 20051
rect 208367 20023 208401 20051
rect 208429 20023 208464 20051
rect 208304 19989 208464 20023
rect 208304 19961 208339 19989
rect 208367 19961 208401 19989
rect 208429 19961 208464 19989
rect 208304 19944 208464 19961
rect 223664 20175 223824 20192
rect 223664 20147 223699 20175
rect 223727 20147 223761 20175
rect 223789 20147 223824 20175
rect 223664 20113 223824 20147
rect 223664 20085 223699 20113
rect 223727 20085 223761 20113
rect 223789 20085 223824 20113
rect 223664 20051 223824 20085
rect 223664 20023 223699 20051
rect 223727 20023 223761 20051
rect 223789 20023 223824 20051
rect 223664 19989 223824 20023
rect 223664 19961 223699 19989
rect 223727 19961 223761 19989
rect 223789 19961 223824 19989
rect 223664 19944 223824 19961
rect 239024 20175 239184 20192
rect 239024 20147 239059 20175
rect 239087 20147 239121 20175
rect 239149 20147 239184 20175
rect 239024 20113 239184 20147
rect 239024 20085 239059 20113
rect 239087 20085 239121 20113
rect 239149 20085 239184 20113
rect 239024 20051 239184 20085
rect 239024 20023 239059 20051
rect 239087 20023 239121 20051
rect 239149 20023 239184 20051
rect 239024 19989 239184 20023
rect 239024 19961 239059 19989
rect 239087 19961 239121 19989
rect 239149 19961 239184 19989
rect 239024 19944 239184 19961
rect 254384 20175 254544 20192
rect 254384 20147 254419 20175
rect 254447 20147 254481 20175
rect 254509 20147 254544 20175
rect 254384 20113 254544 20147
rect 254384 20085 254419 20113
rect 254447 20085 254481 20113
rect 254509 20085 254544 20113
rect 254384 20051 254544 20085
rect 254384 20023 254419 20051
rect 254447 20023 254481 20051
rect 254509 20023 254544 20051
rect 254384 19989 254544 20023
rect 254384 19961 254419 19989
rect 254447 19961 254481 19989
rect 254509 19961 254544 19989
rect 254384 19944 254544 19961
rect 269744 20175 269904 20192
rect 269744 20147 269779 20175
rect 269807 20147 269841 20175
rect 269869 20147 269904 20175
rect 269744 20113 269904 20147
rect 269744 20085 269779 20113
rect 269807 20085 269841 20113
rect 269869 20085 269904 20113
rect 269744 20051 269904 20085
rect 269744 20023 269779 20051
rect 269807 20023 269841 20051
rect 269869 20023 269904 20051
rect 269744 19989 269904 20023
rect 269744 19961 269779 19989
rect 269807 19961 269841 19989
rect 269869 19961 269904 19989
rect 269744 19944 269904 19961
rect 158169 14147 158217 14175
rect 158245 14147 158279 14175
rect 158307 14147 158341 14175
rect 158369 14147 158403 14175
rect 158431 14147 158479 14175
rect 158169 14113 158479 14147
rect 158169 14085 158217 14113
rect 158245 14085 158279 14113
rect 158307 14085 158341 14113
rect 158369 14085 158403 14113
rect 158431 14085 158479 14113
rect 158169 14051 158479 14085
rect 158169 14023 158217 14051
rect 158245 14023 158279 14051
rect 158307 14023 158341 14051
rect 158369 14023 158403 14051
rect 158431 14023 158479 14051
rect 158169 13989 158479 14023
rect 158169 13961 158217 13989
rect 158245 13961 158279 13989
rect 158307 13961 158341 13989
rect 158369 13961 158403 13989
rect 158431 13961 158479 13989
rect 158169 5175 158479 13961
rect 169904 14175 170064 14192
rect 169904 14147 169939 14175
rect 169967 14147 170001 14175
rect 170029 14147 170064 14175
rect 169904 14113 170064 14147
rect 169904 14085 169939 14113
rect 169967 14085 170001 14113
rect 170029 14085 170064 14113
rect 169904 14051 170064 14085
rect 169904 14023 169939 14051
rect 169967 14023 170001 14051
rect 170029 14023 170064 14051
rect 169904 13989 170064 14023
rect 169904 13961 169939 13989
rect 169967 13961 170001 13989
rect 170029 13961 170064 13989
rect 169904 13944 170064 13961
rect 185264 14175 185424 14192
rect 185264 14147 185299 14175
rect 185327 14147 185361 14175
rect 185389 14147 185424 14175
rect 185264 14113 185424 14147
rect 185264 14085 185299 14113
rect 185327 14085 185361 14113
rect 185389 14085 185424 14113
rect 185264 14051 185424 14085
rect 185264 14023 185299 14051
rect 185327 14023 185361 14051
rect 185389 14023 185424 14051
rect 185264 13989 185424 14023
rect 185264 13961 185299 13989
rect 185327 13961 185361 13989
rect 185389 13961 185424 13989
rect 185264 13944 185424 13961
rect 200624 14175 200784 14192
rect 200624 14147 200659 14175
rect 200687 14147 200721 14175
rect 200749 14147 200784 14175
rect 200624 14113 200784 14147
rect 200624 14085 200659 14113
rect 200687 14085 200721 14113
rect 200749 14085 200784 14113
rect 200624 14051 200784 14085
rect 200624 14023 200659 14051
rect 200687 14023 200721 14051
rect 200749 14023 200784 14051
rect 200624 13989 200784 14023
rect 200624 13961 200659 13989
rect 200687 13961 200721 13989
rect 200749 13961 200784 13989
rect 200624 13944 200784 13961
rect 215984 14175 216144 14192
rect 215984 14147 216019 14175
rect 216047 14147 216081 14175
rect 216109 14147 216144 14175
rect 215984 14113 216144 14147
rect 215984 14085 216019 14113
rect 216047 14085 216081 14113
rect 216109 14085 216144 14113
rect 215984 14051 216144 14085
rect 215984 14023 216019 14051
rect 216047 14023 216081 14051
rect 216109 14023 216144 14051
rect 215984 13989 216144 14023
rect 215984 13961 216019 13989
rect 216047 13961 216081 13989
rect 216109 13961 216144 13989
rect 215984 13944 216144 13961
rect 231344 14175 231504 14192
rect 231344 14147 231379 14175
rect 231407 14147 231441 14175
rect 231469 14147 231504 14175
rect 231344 14113 231504 14147
rect 231344 14085 231379 14113
rect 231407 14085 231441 14113
rect 231469 14085 231504 14113
rect 231344 14051 231504 14085
rect 231344 14023 231379 14051
rect 231407 14023 231441 14051
rect 231469 14023 231504 14051
rect 231344 13989 231504 14023
rect 231344 13961 231379 13989
rect 231407 13961 231441 13989
rect 231469 13961 231504 13989
rect 231344 13944 231504 13961
rect 246704 14175 246864 14192
rect 246704 14147 246739 14175
rect 246767 14147 246801 14175
rect 246829 14147 246864 14175
rect 246704 14113 246864 14147
rect 246704 14085 246739 14113
rect 246767 14085 246801 14113
rect 246829 14085 246864 14113
rect 246704 14051 246864 14085
rect 246704 14023 246739 14051
rect 246767 14023 246801 14051
rect 246829 14023 246864 14051
rect 246704 13989 246864 14023
rect 246704 13961 246739 13989
rect 246767 13961 246801 13989
rect 246829 13961 246864 13989
rect 246704 13944 246864 13961
rect 262064 14175 262224 14192
rect 262064 14147 262099 14175
rect 262127 14147 262161 14175
rect 262189 14147 262224 14175
rect 262064 14113 262224 14147
rect 262064 14085 262099 14113
rect 262127 14085 262161 14113
rect 262189 14085 262224 14113
rect 262064 14051 262224 14085
rect 262064 14023 262099 14051
rect 262127 14023 262161 14051
rect 262189 14023 262224 14051
rect 262064 13989 262224 14023
rect 262064 13961 262099 13989
rect 262127 13961 262161 13989
rect 262189 13961 262224 13989
rect 262064 13944 262224 13961
rect 162224 11175 162384 11192
rect 162224 11147 162259 11175
rect 162287 11147 162321 11175
rect 162349 11147 162384 11175
rect 162224 11113 162384 11147
rect 162224 11085 162259 11113
rect 162287 11085 162321 11113
rect 162349 11085 162384 11113
rect 162224 11051 162384 11085
rect 162224 11023 162259 11051
rect 162287 11023 162321 11051
rect 162349 11023 162384 11051
rect 162224 10989 162384 11023
rect 162224 10961 162259 10989
rect 162287 10961 162321 10989
rect 162349 10961 162384 10989
rect 162224 10944 162384 10961
rect 177584 11175 177744 11192
rect 177584 11147 177619 11175
rect 177647 11147 177681 11175
rect 177709 11147 177744 11175
rect 177584 11113 177744 11147
rect 177584 11085 177619 11113
rect 177647 11085 177681 11113
rect 177709 11085 177744 11113
rect 177584 11051 177744 11085
rect 177584 11023 177619 11051
rect 177647 11023 177681 11051
rect 177709 11023 177744 11051
rect 177584 10989 177744 11023
rect 177584 10961 177619 10989
rect 177647 10961 177681 10989
rect 177709 10961 177744 10989
rect 177584 10944 177744 10961
rect 192944 11175 193104 11192
rect 192944 11147 192979 11175
rect 193007 11147 193041 11175
rect 193069 11147 193104 11175
rect 192944 11113 193104 11147
rect 192944 11085 192979 11113
rect 193007 11085 193041 11113
rect 193069 11085 193104 11113
rect 192944 11051 193104 11085
rect 192944 11023 192979 11051
rect 193007 11023 193041 11051
rect 193069 11023 193104 11051
rect 192944 10989 193104 11023
rect 192944 10961 192979 10989
rect 193007 10961 193041 10989
rect 193069 10961 193104 10989
rect 192944 10944 193104 10961
rect 208304 11175 208464 11192
rect 208304 11147 208339 11175
rect 208367 11147 208401 11175
rect 208429 11147 208464 11175
rect 208304 11113 208464 11147
rect 208304 11085 208339 11113
rect 208367 11085 208401 11113
rect 208429 11085 208464 11113
rect 208304 11051 208464 11085
rect 208304 11023 208339 11051
rect 208367 11023 208401 11051
rect 208429 11023 208464 11051
rect 208304 10989 208464 11023
rect 208304 10961 208339 10989
rect 208367 10961 208401 10989
rect 208429 10961 208464 10989
rect 208304 10944 208464 10961
rect 223664 11175 223824 11192
rect 223664 11147 223699 11175
rect 223727 11147 223761 11175
rect 223789 11147 223824 11175
rect 223664 11113 223824 11147
rect 223664 11085 223699 11113
rect 223727 11085 223761 11113
rect 223789 11085 223824 11113
rect 223664 11051 223824 11085
rect 223664 11023 223699 11051
rect 223727 11023 223761 11051
rect 223789 11023 223824 11051
rect 223664 10989 223824 11023
rect 223664 10961 223699 10989
rect 223727 10961 223761 10989
rect 223789 10961 223824 10989
rect 223664 10944 223824 10961
rect 239024 11175 239184 11192
rect 239024 11147 239059 11175
rect 239087 11147 239121 11175
rect 239149 11147 239184 11175
rect 239024 11113 239184 11147
rect 239024 11085 239059 11113
rect 239087 11085 239121 11113
rect 239149 11085 239184 11113
rect 239024 11051 239184 11085
rect 239024 11023 239059 11051
rect 239087 11023 239121 11051
rect 239149 11023 239184 11051
rect 239024 10989 239184 11023
rect 239024 10961 239059 10989
rect 239087 10961 239121 10989
rect 239149 10961 239184 10989
rect 239024 10944 239184 10961
rect 254384 11175 254544 11192
rect 254384 11147 254419 11175
rect 254447 11147 254481 11175
rect 254509 11147 254544 11175
rect 254384 11113 254544 11147
rect 254384 11085 254419 11113
rect 254447 11085 254481 11113
rect 254509 11085 254544 11113
rect 254384 11051 254544 11085
rect 254384 11023 254419 11051
rect 254447 11023 254481 11051
rect 254509 11023 254544 11051
rect 254384 10989 254544 11023
rect 254384 10961 254419 10989
rect 254447 10961 254481 10989
rect 254509 10961 254544 10989
rect 254384 10944 254544 10961
rect 269744 11175 269904 11192
rect 269744 11147 269779 11175
rect 269807 11147 269841 11175
rect 269869 11147 269904 11175
rect 269744 11113 269904 11147
rect 269744 11085 269779 11113
rect 269807 11085 269841 11113
rect 269869 11085 269904 11113
rect 269744 11051 269904 11085
rect 269744 11023 269779 11051
rect 269807 11023 269841 11051
rect 269869 11023 269904 11051
rect 269744 10989 269904 11023
rect 269744 10961 269779 10989
rect 269807 10961 269841 10989
rect 269869 10961 269904 10989
rect 269744 10944 269904 10961
rect 158169 5147 158217 5175
rect 158245 5147 158279 5175
rect 158307 5147 158341 5175
rect 158369 5147 158403 5175
rect 158431 5147 158479 5175
rect 158169 5113 158479 5147
rect 158169 5085 158217 5113
rect 158245 5085 158279 5113
rect 158307 5085 158341 5113
rect 158369 5085 158403 5113
rect 158431 5085 158479 5113
rect 158169 5051 158479 5085
rect 158169 5023 158217 5051
rect 158245 5023 158279 5051
rect 158307 5023 158341 5051
rect 158369 5023 158403 5051
rect 158431 5023 158479 5051
rect 158169 4989 158479 5023
rect 158169 4961 158217 4989
rect 158245 4961 158279 4989
rect 158307 4961 158341 4989
rect 158369 4961 158403 4989
rect 158431 4961 158479 4989
rect 158169 -560 158479 4961
rect 158169 -588 158217 -560
rect 158245 -588 158279 -560
rect 158307 -588 158341 -560
rect 158369 -588 158403 -560
rect 158431 -588 158479 -560
rect 158169 -622 158479 -588
rect 158169 -650 158217 -622
rect 158245 -650 158279 -622
rect 158307 -650 158341 -622
rect 158369 -650 158403 -622
rect 158431 -650 158479 -622
rect 158169 -684 158479 -650
rect 158169 -712 158217 -684
rect 158245 -712 158279 -684
rect 158307 -712 158341 -684
rect 158369 -712 158403 -684
rect 158431 -712 158479 -684
rect 158169 -746 158479 -712
rect 158169 -774 158217 -746
rect 158245 -774 158279 -746
rect 158307 -774 158341 -746
rect 158369 -774 158403 -746
rect 158431 -774 158479 -746
rect 158169 -822 158479 -774
rect 171669 2175 171979 6401
rect 171669 2147 171717 2175
rect 171745 2147 171779 2175
rect 171807 2147 171841 2175
rect 171869 2147 171903 2175
rect 171931 2147 171979 2175
rect 171669 2113 171979 2147
rect 171669 2085 171717 2113
rect 171745 2085 171779 2113
rect 171807 2085 171841 2113
rect 171869 2085 171903 2113
rect 171931 2085 171979 2113
rect 171669 2051 171979 2085
rect 171669 2023 171717 2051
rect 171745 2023 171779 2051
rect 171807 2023 171841 2051
rect 171869 2023 171903 2051
rect 171931 2023 171979 2051
rect 171669 1989 171979 2023
rect 171669 1961 171717 1989
rect 171745 1961 171779 1989
rect 171807 1961 171841 1989
rect 171869 1961 171903 1989
rect 171931 1961 171979 1989
rect 171669 -80 171979 1961
rect 171669 -108 171717 -80
rect 171745 -108 171779 -80
rect 171807 -108 171841 -80
rect 171869 -108 171903 -80
rect 171931 -108 171979 -80
rect 171669 -142 171979 -108
rect 171669 -170 171717 -142
rect 171745 -170 171779 -142
rect 171807 -170 171841 -142
rect 171869 -170 171903 -142
rect 171931 -170 171979 -142
rect 171669 -204 171979 -170
rect 171669 -232 171717 -204
rect 171745 -232 171779 -204
rect 171807 -232 171841 -204
rect 171869 -232 171903 -204
rect 171931 -232 171979 -204
rect 171669 -266 171979 -232
rect 171669 -294 171717 -266
rect 171745 -294 171779 -266
rect 171807 -294 171841 -266
rect 171869 -294 171903 -266
rect 171931 -294 171979 -266
rect 171669 -822 171979 -294
rect 173529 5175 173839 6401
rect 173529 5147 173577 5175
rect 173605 5147 173639 5175
rect 173667 5147 173701 5175
rect 173729 5147 173763 5175
rect 173791 5147 173839 5175
rect 173529 5113 173839 5147
rect 173529 5085 173577 5113
rect 173605 5085 173639 5113
rect 173667 5085 173701 5113
rect 173729 5085 173763 5113
rect 173791 5085 173839 5113
rect 173529 5051 173839 5085
rect 173529 5023 173577 5051
rect 173605 5023 173639 5051
rect 173667 5023 173701 5051
rect 173729 5023 173763 5051
rect 173791 5023 173839 5051
rect 173529 4989 173839 5023
rect 173529 4961 173577 4989
rect 173605 4961 173639 4989
rect 173667 4961 173701 4989
rect 173729 4961 173763 4989
rect 173791 4961 173839 4989
rect 173529 -560 173839 4961
rect 173529 -588 173577 -560
rect 173605 -588 173639 -560
rect 173667 -588 173701 -560
rect 173729 -588 173763 -560
rect 173791 -588 173839 -560
rect 173529 -622 173839 -588
rect 173529 -650 173577 -622
rect 173605 -650 173639 -622
rect 173667 -650 173701 -622
rect 173729 -650 173763 -622
rect 173791 -650 173839 -622
rect 173529 -684 173839 -650
rect 173529 -712 173577 -684
rect 173605 -712 173639 -684
rect 173667 -712 173701 -684
rect 173729 -712 173763 -684
rect 173791 -712 173839 -684
rect 173529 -746 173839 -712
rect 173529 -774 173577 -746
rect 173605 -774 173639 -746
rect 173667 -774 173701 -746
rect 173729 -774 173763 -746
rect 173791 -774 173839 -746
rect 173529 -822 173839 -774
rect 187029 2175 187339 6401
rect 187029 2147 187077 2175
rect 187105 2147 187139 2175
rect 187167 2147 187201 2175
rect 187229 2147 187263 2175
rect 187291 2147 187339 2175
rect 187029 2113 187339 2147
rect 187029 2085 187077 2113
rect 187105 2085 187139 2113
rect 187167 2085 187201 2113
rect 187229 2085 187263 2113
rect 187291 2085 187339 2113
rect 187029 2051 187339 2085
rect 187029 2023 187077 2051
rect 187105 2023 187139 2051
rect 187167 2023 187201 2051
rect 187229 2023 187263 2051
rect 187291 2023 187339 2051
rect 187029 1989 187339 2023
rect 187029 1961 187077 1989
rect 187105 1961 187139 1989
rect 187167 1961 187201 1989
rect 187229 1961 187263 1989
rect 187291 1961 187339 1989
rect 187029 -80 187339 1961
rect 187029 -108 187077 -80
rect 187105 -108 187139 -80
rect 187167 -108 187201 -80
rect 187229 -108 187263 -80
rect 187291 -108 187339 -80
rect 187029 -142 187339 -108
rect 187029 -170 187077 -142
rect 187105 -170 187139 -142
rect 187167 -170 187201 -142
rect 187229 -170 187263 -142
rect 187291 -170 187339 -142
rect 187029 -204 187339 -170
rect 187029 -232 187077 -204
rect 187105 -232 187139 -204
rect 187167 -232 187201 -204
rect 187229 -232 187263 -204
rect 187291 -232 187339 -204
rect 187029 -266 187339 -232
rect 187029 -294 187077 -266
rect 187105 -294 187139 -266
rect 187167 -294 187201 -266
rect 187229 -294 187263 -266
rect 187291 -294 187339 -266
rect 187029 -822 187339 -294
rect 188889 5175 189199 6401
rect 188889 5147 188937 5175
rect 188965 5147 188999 5175
rect 189027 5147 189061 5175
rect 189089 5147 189123 5175
rect 189151 5147 189199 5175
rect 188889 5113 189199 5147
rect 188889 5085 188937 5113
rect 188965 5085 188999 5113
rect 189027 5085 189061 5113
rect 189089 5085 189123 5113
rect 189151 5085 189199 5113
rect 188889 5051 189199 5085
rect 188889 5023 188937 5051
rect 188965 5023 188999 5051
rect 189027 5023 189061 5051
rect 189089 5023 189123 5051
rect 189151 5023 189199 5051
rect 188889 4989 189199 5023
rect 188889 4961 188937 4989
rect 188965 4961 188999 4989
rect 189027 4961 189061 4989
rect 189089 4961 189123 4989
rect 189151 4961 189199 4989
rect 188889 -560 189199 4961
rect 188889 -588 188937 -560
rect 188965 -588 188999 -560
rect 189027 -588 189061 -560
rect 189089 -588 189123 -560
rect 189151 -588 189199 -560
rect 188889 -622 189199 -588
rect 188889 -650 188937 -622
rect 188965 -650 188999 -622
rect 189027 -650 189061 -622
rect 189089 -650 189123 -622
rect 189151 -650 189199 -622
rect 188889 -684 189199 -650
rect 188889 -712 188937 -684
rect 188965 -712 188999 -684
rect 189027 -712 189061 -684
rect 189089 -712 189123 -684
rect 189151 -712 189199 -684
rect 188889 -746 189199 -712
rect 188889 -774 188937 -746
rect 188965 -774 188999 -746
rect 189027 -774 189061 -746
rect 189089 -774 189123 -746
rect 189151 -774 189199 -746
rect 188889 -822 189199 -774
rect 202389 2175 202699 6401
rect 202389 2147 202437 2175
rect 202465 2147 202499 2175
rect 202527 2147 202561 2175
rect 202589 2147 202623 2175
rect 202651 2147 202699 2175
rect 202389 2113 202699 2147
rect 202389 2085 202437 2113
rect 202465 2085 202499 2113
rect 202527 2085 202561 2113
rect 202589 2085 202623 2113
rect 202651 2085 202699 2113
rect 202389 2051 202699 2085
rect 202389 2023 202437 2051
rect 202465 2023 202499 2051
rect 202527 2023 202561 2051
rect 202589 2023 202623 2051
rect 202651 2023 202699 2051
rect 202389 1989 202699 2023
rect 202389 1961 202437 1989
rect 202465 1961 202499 1989
rect 202527 1961 202561 1989
rect 202589 1961 202623 1989
rect 202651 1961 202699 1989
rect 202389 -80 202699 1961
rect 202389 -108 202437 -80
rect 202465 -108 202499 -80
rect 202527 -108 202561 -80
rect 202589 -108 202623 -80
rect 202651 -108 202699 -80
rect 202389 -142 202699 -108
rect 202389 -170 202437 -142
rect 202465 -170 202499 -142
rect 202527 -170 202561 -142
rect 202589 -170 202623 -142
rect 202651 -170 202699 -142
rect 202389 -204 202699 -170
rect 202389 -232 202437 -204
rect 202465 -232 202499 -204
rect 202527 -232 202561 -204
rect 202589 -232 202623 -204
rect 202651 -232 202699 -204
rect 202389 -266 202699 -232
rect 202389 -294 202437 -266
rect 202465 -294 202499 -266
rect 202527 -294 202561 -266
rect 202589 -294 202623 -266
rect 202651 -294 202699 -266
rect 202389 -822 202699 -294
rect 204249 5175 204559 6401
rect 204249 5147 204297 5175
rect 204325 5147 204359 5175
rect 204387 5147 204421 5175
rect 204449 5147 204483 5175
rect 204511 5147 204559 5175
rect 204249 5113 204559 5147
rect 204249 5085 204297 5113
rect 204325 5085 204359 5113
rect 204387 5085 204421 5113
rect 204449 5085 204483 5113
rect 204511 5085 204559 5113
rect 204249 5051 204559 5085
rect 204249 5023 204297 5051
rect 204325 5023 204359 5051
rect 204387 5023 204421 5051
rect 204449 5023 204483 5051
rect 204511 5023 204559 5051
rect 204249 4989 204559 5023
rect 204249 4961 204297 4989
rect 204325 4961 204359 4989
rect 204387 4961 204421 4989
rect 204449 4961 204483 4989
rect 204511 4961 204559 4989
rect 204249 -560 204559 4961
rect 204249 -588 204297 -560
rect 204325 -588 204359 -560
rect 204387 -588 204421 -560
rect 204449 -588 204483 -560
rect 204511 -588 204559 -560
rect 204249 -622 204559 -588
rect 204249 -650 204297 -622
rect 204325 -650 204359 -622
rect 204387 -650 204421 -622
rect 204449 -650 204483 -622
rect 204511 -650 204559 -622
rect 204249 -684 204559 -650
rect 204249 -712 204297 -684
rect 204325 -712 204359 -684
rect 204387 -712 204421 -684
rect 204449 -712 204483 -684
rect 204511 -712 204559 -684
rect 204249 -746 204559 -712
rect 204249 -774 204297 -746
rect 204325 -774 204359 -746
rect 204387 -774 204421 -746
rect 204449 -774 204483 -746
rect 204511 -774 204559 -746
rect 204249 -822 204559 -774
rect 217749 2175 218059 6401
rect 217749 2147 217797 2175
rect 217825 2147 217859 2175
rect 217887 2147 217921 2175
rect 217949 2147 217983 2175
rect 218011 2147 218059 2175
rect 217749 2113 218059 2147
rect 217749 2085 217797 2113
rect 217825 2085 217859 2113
rect 217887 2085 217921 2113
rect 217949 2085 217983 2113
rect 218011 2085 218059 2113
rect 217749 2051 218059 2085
rect 217749 2023 217797 2051
rect 217825 2023 217859 2051
rect 217887 2023 217921 2051
rect 217949 2023 217983 2051
rect 218011 2023 218059 2051
rect 217749 1989 218059 2023
rect 217749 1961 217797 1989
rect 217825 1961 217859 1989
rect 217887 1961 217921 1989
rect 217949 1961 217983 1989
rect 218011 1961 218059 1989
rect 217749 -80 218059 1961
rect 217749 -108 217797 -80
rect 217825 -108 217859 -80
rect 217887 -108 217921 -80
rect 217949 -108 217983 -80
rect 218011 -108 218059 -80
rect 217749 -142 218059 -108
rect 217749 -170 217797 -142
rect 217825 -170 217859 -142
rect 217887 -170 217921 -142
rect 217949 -170 217983 -142
rect 218011 -170 218059 -142
rect 217749 -204 218059 -170
rect 217749 -232 217797 -204
rect 217825 -232 217859 -204
rect 217887 -232 217921 -204
rect 217949 -232 217983 -204
rect 218011 -232 218059 -204
rect 217749 -266 218059 -232
rect 217749 -294 217797 -266
rect 217825 -294 217859 -266
rect 217887 -294 217921 -266
rect 217949 -294 217983 -266
rect 218011 -294 218059 -266
rect 217749 -822 218059 -294
rect 219609 5175 219919 6401
rect 219609 5147 219657 5175
rect 219685 5147 219719 5175
rect 219747 5147 219781 5175
rect 219809 5147 219843 5175
rect 219871 5147 219919 5175
rect 219609 5113 219919 5147
rect 219609 5085 219657 5113
rect 219685 5085 219719 5113
rect 219747 5085 219781 5113
rect 219809 5085 219843 5113
rect 219871 5085 219919 5113
rect 219609 5051 219919 5085
rect 219609 5023 219657 5051
rect 219685 5023 219719 5051
rect 219747 5023 219781 5051
rect 219809 5023 219843 5051
rect 219871 5023 219919 5051
rect 219609 4989 219919 5023
rect 219609 4961 219657 4989
rect 219685 4961 219719 4989
rect 219747 4961 219781 4989
rect 219809 4961 219843 4989
rect 219871 4961 219919 4989
rect 219609 -560 219919 4961
rect 219609 -588 219657 -560
rect 219685 -588 219719 -560
rect 219747 -588 219781 -560
rect 219809 -588 219843 -560
rect 219871 -588 219919 -560
rect 219609 -622 219919 -588
rect 219609 -650 219657 -622
rect 219685 -650 219719 -622
rect 219747 -650 219781 -622
rect 219809 -650 219843 -622
rect 219871 -650 219919 -622
rect 219609 -684 219919 -650
rect 219609 -712 219657 -684
rect 219685 -712 219719 -684
rect 219747 -712 219781 -684
rect 219809 -712 219843 -684
rect 219871 -712 219919 -684
rect 219609 -746 219919 -712
rect 219609 -774 219657 -746
rect 219685 -774 219719 -746
rect 219747 -774 219781 -746
rect 219809 -774 219843 -746
rect 219871 -774 219919 -746
rect 219609 -822 219919 -774
rect 233109 2175 233419 6401
rect 233109 2147 233157 2175
rect 233185 2147 233219 2175
rect 233247 2147 233281 2175
rect 233309 2147 233343 2175
rect 233371 2147 233419 2175
rect 233109 2113 233419 2147
rect 233109 2085 233157 2113
rect 233185 2085 233219 2113
rect 233247 2085 233281 2113
rect 233309 2085 233343 2113
rect 233371 2085 233419 2113
rect 233109 2051 233419 2085
rect 233109 2023 233157 2051
rect 233185 2023 233219 2051
rect 233247 2023 233281 2051
rect 233309 2023 233343 2051
rect 233371 2023 233419 2051
rect 233109 1989 233419 2023
rect 233109 1961 233157 1989
rect 233185 1961 233219 1989
rect 233247 1961 233281 1989
rect 233309 1961 233343 1989
rect 233371 1961 233419 1989
rect 233109 -80 233419 1961
rect 233109 -108 233157 -80
rect 233185 -108 233219 -80
rect 233247 -108 233281 -80
rect 233309 -108 233343 -80
rect 233371 -108 233419 -80
rect 233109 -142 233419 -108
rect 233109 -170 233157 -142
rect 233185 -170 233219 -142
rect 233247 -170 233281 -142
rect 233309 -170 233343 -142
rect 233371 -170 233419 -142
rect 233109 -204 233419 -170
rect 233109 -232 233157 -204
rect 233185 -232 233219 -204
rect 233247 -232 233281 -204
rect 233309 -232 233343 -204
rect 233371 -232 233419 -204
rect 233109 -266 233419 -232
rect 233109 -294 233157 -266
rect 233185 -294 233219 -266
rect 233247 -294 233281 -266
rect 233309 -294 233343 -266
rect 233371 -294 233419 -266
rect 233109 -822 233419 -294
rect 234969 5175 235279 6401
rect 234969 5147 235017 5175
rect 235045 5147 235079 5175
rect 235107 5147 235141 5175
rect 235169 5147 235203 5175
rect 235231 5147 235279 5175
rect 234969 5113 235279 5147
rect 234969 5085 235017 5113
rect 235045 5085 235079 5113
rect 235107 5085 235141 5113
rect 235169 5085 235203 5113
rect 235231 5085 235279 5113
rect 234969 5051 235279 5085
rect 234969 5023 235017 5051
rect 235045 5023 235079 5051
rect 235107 5023 235141 5051
rect 235169 5023 235203 5051
rect 235231 5023 235279 5051
rect 234969 4989 235279 5023
rect 234969 4961 235017 4989
rect 235045 4961 235079 4989
rect 235107 4961 235141 4989
rect 235169 4961 235203 4989
rect 235231 4961 235279 4989
rect 234969 -560 235279 4961
rect 234969 -588 235017 -560
rect 235045 -588 235079 -560
rect 235107 -588 235141 -560
rect 235169 -588 235203 -560
rect 235231 -588 235279 -560
rect 234969 -622 235279 -588
rect 234969 -650 235017 -622
rect 235045 -650 235079 -622
rect 235107 -650 235141 -622
rect 235169 -650 235203 -622
rect 235231 -650 235279 -622
rect 234969 -684 235279 -650
rect 234969 -712 235017 -684
rect 235045 -712 235079 -684
rect 235107 -712 235141 -684
rect 235169 -712 235203 -684
rect 235231 -712 235279 -684
rect 234969 -746 235279 -712
rect 234969 -774 235017 -746
rect 235045 -774 235079 -746
rect 235107 -774 235141 -746
rect 235169 -774 235203 -746
rect 235231 -774 235279 -746
rect 234969 -822 235279 -774
rect 248469 2175 248779 6401
rect 248469 2147 248517 2175
rect 248545 2147 248579 2175
rect 248607 2147 248641 2175
rect 248669 2147 248703 2175
rect 248731 2147 248779 2175
rect 248469 2113 248779 2147
rect 248469 2085 248517 2113
rect 248545 2085 248579 2113
rect 248607 2085 248641 2113
rect 248669 2085 248703 2113
rect 248731 2085 248779 2113
rect 248469 2051 248779 2085
rect 248469 2023 248517 2051
rect 248545 2023 248579 2051
rect 248607 2023 248641 2051
rect 248669 2023 248703 2051
rect 248731 2023 248779 2051
rect 248469 1989 248779 2023
rect 248469 1961 248517 1989
rect 248545 1961 248579 1989
rect 248607 1961 248641 1989
rect 248669 1961 248703 1989
rect 248731 1961 248779 1989
rect 248469 -80 248779 1961
rect 248469 -108 248517 -80
rect 248545 -108 248579 -80
rect 248607 -108 248641 -80
rect 248669 -108 248703 -80
rect 248731 -108 248779 -80
rect 248469 -142 248779 -108
rect 248469 -170 248517 -142
rect 248545 -170 248579 -142
rect 248607 -170 248641 -142
rect 248669 -170 248703 -142
rect 248731 -170 248779 -142
rect 248469 -204 248779 -170
rect 248469 -232 248517 -204
rect 248545 -232 248579 -204
rect 248607 -232 248641 -204
rect 248669 -232 248703 -204
rect 248731 -232 248779 -204
rect 248469 -266 248779 -232
rect 248469 -294 248517 -266
rect 248545 -294 248579 -266
rect 248607 -294 248641 -266
rect 248669 -294 248703 -266
rect 248731 -294 248779 -266
rect 248469 -822 248779 -294
rect 250329 5175 250639 6401
rect 250329 5147 250377 5175
rect 250405 5147 250439 5175
rect 250467 5147 250501 5175
rect 250529 5147 250563 5175
rect 250591 5147 250639 5175
rect 250329 5113 250639 5147
rect 250329 5085 250377 5113
rect 250405 5085 250439 5113
rect 250467 5085 250501 5113
rect 250529 5085 250563 5113
rect 250591 5085 250639 5113
rect 250329 5051 250639 5085
rect 250329 5023 250377 5051
rect 250405 5023 250439 5051
rect 250467 5023 250501 5051
rect 250529 5023 250563 5051
rect 250591 5023 250639 5051
rect 250329 4989 250639 5023
rect 250329 4961 250377 4989
rect 250405 4961 250439 4989
rect 250467 4961 250501 4989
rect 250529 4961 250563 4989
rect 250591 4961 250639 4989
rect 250329 -560 250639 4961
rect 250329 -588 250377 -560
rect 250405 -588 250439 -560
rect 250467 -588 250501 -560
rect 250529 -588 250563 -560
rect 250591 -588 250639 -560
rect 250329 -622 250639 -588
rect 250329 -650 250377 -622
rect 250405 -650 250439 -622
rect 250467 -650 250501 -622
rect 250529 -650 250563 -622
rect 250591 -650 250639 -622
rect 250329 -684 250639 -650
rect 250329 -712 250377 -684
rect 250405 -712 250439 -684
rect 250467 -712 250501 -684
rect 250529 -712 250563 -684
rect 250591 -712 250639 -684
rect 250329 -746 250639 -712
rect 250329 -774 250377 -746
rect 250405 -774 250439 -746
rect 250467 -774 250501 -746
rect 250529 -774 250563 -746
rect 250591 -774 250639 -746
rect 250329 -822 250639 -774
rect 263829 2175 264139 6401
rect 263829 2147 263877 2175
rect 263905 2147 263939 2175
rect 263967 2147 264001 2175
rect 264029 2147 264063 2175
rect 264091 2147 264139 2175
rect 263829 2113 264139 2147
rect 263829 2085 263877 2113
rect 263905 2085 263939 2113
rect 263967 2085 264001 2113
rect 264029 2085 264063 2113
rect 264091 2085 264139 2113
rect 263829 2051 264139 2085
rect 263829 2023 263877 2051
rect 263905 2023 263939 2051
rect 263967 2023 264001 2051
rect 264029 2023 264063 2051
rect 264091 2023 264139 2051
rect 263829 1989 264139 2023
rect 263829 1961 263877 1989
rect 263905 1961 263939 1989
rect 263967 1961 264001 1989
rect 264029 1961 264063 1989
rect 264091 1961 264139 1989
rect 263829 -80 264139 1961
rect 263829 -108 263877 -80
rect 263905 -108 263939 -80
rect 263967 -108 264001 -80
rect 264029 -108 264063 -80
rect 264091 -108 264139 -80
rect 263829 -142 264139 -108
rect 263829 -170 263877 -142
rect 263905 -170 263939 -142
rect 263967 -170 264001 -142
rect 264029 -170 264063 -142
rect 264091 -170 264139 -142
rect 263829 -204 264139 -170
rect 263829 -232 263877 -204
rect 263905 -232 263939 -204
rect 263967 -232 264001 -204
rect 264029 -232 264063 -204
rect 264091 -232 264139 -204
rect 263829 -266 264139 -232
rect 263829 -294 263877 -266
rect 263905 -294 263939 -266
rect 263967 -294 264001 -266
rect 264029 -294 264063 -266
rect 264091 -294 264139 -266
rect 263829 -822 264139 -294
rect 265689 5175 265999 6401
rect 265689 5147 265737 5175
rect 265765 5147 265799 5175
rect 265827 5147 265861 5175
rect 265889 5147 265923 5175
rect 265951 5147 265999 5175
rect 265689 5113 265999 5147
rect 265689 5085 265737 5113
rect 265765 5085 265799 5113
rect 265827 5085 265861 5113
rect 265889 5085 265923 5113
rect 265951 5085 265999 5113
rect 265689 5051 265999 5085
rect 265689 5023 265737 5051
rect 265765 5023 265799 5051
rect 265827 5023 265861 5051
rect 265889 5023 265923 5051
rect 265951 5023 265999 5051
rect 265689 4989 265999 5023
rect 265689 4961 265737 4989
rect 265765 4961 265799 4989
rect 265827 4961 265861 4989
rect 265889 4961 265923 4989
rect 265951 4961 265999 4989
rect 265689 -560 265999 4961
rect 275926 3570 275954 137942
rect 275982 16842 276010 138838
rect 276038 43218 276066 140630
rect 276038 43185 276066 43190
rect 276094 139314 276122 139319
rect 276094 23394 276122 139286
rect 276150 63042 276178 141974
rect 276822 141554 276850 141559
rect 276150 63009 276178 63014
rect 276766 140210 276794 140215
rect 276766 36610 276794 140182
rect 276822 56434 276850 141526
rect 276878 82866 276906 143318
rect 276934 102690 276962 144662
rect 276990 122514 277018 146006
rect 276990 122481 277018 122486
rect 279189 146023 279237 146051
rect 279265 146023 279299 146051
rect 279327 146023 279361 146051
rect 279389 146023 279423 146051
rect 279451 146023 279499 146051
rect 279189 145989 279499 146023
rect 279189 145961 279237 145989
rect 279265 145961 279299 145989
rect 279327 145961 279361 145989
rect 279389 145961 279423 145989
rect 279451 145961 279499 145989
rect 279189 137175 279499 145961
rect 279189 137147 279237 137175
rect 279265 137147 279299 137175
rect 279327 137147 279361 137175
rect 279389 137147 279423 137175
rect 279451 137147 279499 137175
rect 279189 137113 279499 137147
rect 279189 137085 279237 137113
rect 279265 137085 279299 137113
rect 279327 137085 279361 137113
rect 279389 137085 279423 137113
rect 279451 137085 279499 137113
rect 279189 137051 279499 137085
rect 279189 137023 279237 137051
rect 279265 137023 279299 137051
rect 279327 137023 279361 137051
rect 279389 137023 279423 137051
rect 279451 137023 279499 137051
rect 279189 136989 279499 137023
rect 279189 136961 279237 136989
rect 279265 136961 279299 136989
rect 279327 136961 279361 136989
rect 279389 136961 279423 136989
rect 279451 136961 279499 136989
rect 279189 128175 279499 136961
rect 279189 128147 279237 128175
rect 279265 128147 279299 128175
rect 279327 128147 279361 128175
rect 279389 128147 279423 128175
rect 279451 128147 279499 128175
rect 279189 128113 279499 128147
rect 279189 128085 279237 128113
rect 279265 128085 279299 128113
rect 279327 128085 279361 128113
rect 279389 128085 279423 128113
rect 279451 128085 279499 128113
rect 279189 128051 279499 128085
rect 279189 128023 279237 128051
rect 279265 128023 279299 128051
rect 279327 128023 279361 128051
rect 279389 128023 279423 128051
rect 279451 128023 279499 128051
rect 279189 127989 279499 128023
rect 279189 127961 279237 127989
rect 279265 127961 279299 127989
rect 279327 127961 279361 127989
rect 279389 127961 279423 127989
rect 279451 127961 279499 127989
rect 276934 102657 276962 102662
rect 279189 119175 279499 127961
rect 279189 119147 279237 119175
rect 279265 119147 279299 119175
rect 279327 119147 279361 119175
rect 279389 119147 279423 119175
rect 279451 119147 279499 119175
rect 279189 119113 279499 119147
rect 279189 119085 279237 119113
rect 279265 119085 279299 119113
rect 279327 119085 279361 119113
rect 279389 119085 279423 119113
rect 279451 119085 279499 119113
rect 279189 119051 279499 119085
rect 279189 119023 279237 119051
rect 279265 119023 279299 119051
rect 279327 119023 279361 119051
rect 279389 119023 279423 119051
rect 279451 119023 279499 119051
rect 279189 118989 279499 119023
rect 279189 118961 279237 118989
rect 279265 118961 279299 118989
rect 279327 118961 279361 118989
rect 279389 118961 279423 118989
rect 279451 118961 279499 118989
rect 279189 110175 279499 118961
rect 279189 110147 279237 110175
rect 279265 110147 279299 110175
rect 279327 110147 279361 110175
rect 279389 110147 279423 110175
rect 279451 110147 279499 110175
rect 279189 110113 279499 110147
rect 279189 110085 279237 110113
rect 279265 110085 279299 110113
rect 279327 110085 279361 110113
rect 279389 110085 279423 110113
rect 279451 110085 279499 110113
rect 279189 110051 279499 110085
rect 279189 110023 279237 110051
rect 279265 110023 279299 110051
rect 279327 110023 279361 110051
rect 279389 110023 279423 110051
rect 279451 110023 279499 110051
rect 279189 109989 279499 110023
rect 279189 109961 279237 109989
rect 279265 109961 279299 109989
rect 279327 109961 279361 109989
rect 279389 109961 279423 109989
rect 279451 109961 279499 109989
rect 276878 82833 276906 82838
rect 279189 101175 279499 109961
rect 279189 101147 279237 101175
rect 279265 101147 279299 101175
rect 279327 101147 279361 101175
rect 279389 101147 279423 101175
rect 279451 101147 279499 101175
rect 279189 101113 279499 101147
rect 279189 101085 279237 101113
rect 279265 101085 279299 101113
rect 279327 101085 279361 101113
rect 279389 101085 279423 101113
rect 279451 101085 279499 101113
rect 279189 101051 279499 101085
rect 279189 101023 279237 101051
rect 279265 101023 279299 101051
rect 279327 101023 279361 101051
rect 279389 101023 279423 101051
rect 279451 101023 279499 101051
rect 279189 100989 279499 101023
rect 279189 100961 279237 100989
rect 279265 100961 279299 100989
rect 279327 100961 279361 100989
rect 279389 100961 279423 100989
rect 279451 100961 279499 100989
rect 279189 92175 279499 100961
rect 279189 92147 279237 92175
rect 279265 92147 279299 92175
rect 279327 92147 279361 92175
rect 279389 92147 279423 92175
rect 279451 92147 279499 92175
rect 279189 92113 279499 92147
rect 279189 92085 279237 92113
rect 279265 92085 279299 92113
rect 279327 92085 279361 92113
rect 279389 92085 279423 92113
rect 279451 92085 279499 92113
rect 279189 92051 279499 92085
rect 279189 92023 279237 92051
rect 279265 92023 279299 92051
rect 279327 92023 279361 92051
rect 279389 92023 279423 92051
rect 279451 92023 279499 92051
rect 279189 91989 279499 92023
rect 279189 91961 279237 91989
rect 279265 91961 279299 91989
rect 279327 91961 279361 91989
rect 279389 91961 279423 91989
rect 279451 91961 279499 91989
rect 279189 83175 279499 91961
rect 279189 83147 279237 83175
rect 279265 83147 279299 83175
rect 279327 83147 279361 83175
rect 279389 83147 279423 83175
rect 279451 83147 279499 83175
rect 279189 83113 279499 83147
rect 279189 83085 279237 83113
rect 279265 83085 279299 83113
rect 279327 83085 279361 83113
rect 279389 83085 279423 83113
rect 279451 83085 279499 83113
rect 279189 83051 279499 83085
rect 279189 83023 279237 83051
rect 279265 83023 279299 83051
rect 279327 83023 279361 83051
rect 279389 83023 279423 83051
rect 279451 83023 279499 83051
rect 279189 82989 279499 83023
rect 279189 82961 279237 82989
rect 279265 82961 279299 82989
rect 279327 82961 279361 82989
rect 279389 82961 279423 82989
rect 279451 82961 279499 82989
rect 276822 56401 276850 56406
rect 279189 74175 279499 82961
rect 279189 74147 279237 74175
rect 279265 74147 279299 74175
rect 279327 74147 279361 74175
rect 279389 74147 279423 74175
rect 279451 74147 279499 74175
rect 279189 74113 279499 74147
rect 279189 74085 279237 74113
rect 279265 74085 279299 74113
rect 279327 74085 279361 74113
rect 279389 74085 279423 74113
rect 279451 74085 279499 74113
rect 279189 74051 279499 74085
rect 279189 74023 279237 74051
rect 279265 74023 279299 74051
rect 279327 74023 279361 74051
rect 279389 74023 279423 74051
rect 279451 74023 279499 74051
rect 279189 73989 279499 74023
rect 279189 73961 279237 73989
rect 279265 73961 279299 73989
rect 279327 73961 279361 73989
rect 279389 73961 279423 73989
rect 279451 73961 279499 73989
rect 279189 65175 279499 73961
rect 279189 65147 279237 65175
rect 279265 65147 279299 65175
rect 279327 65147 279361 65175
rect 279389 65147 279423 65175
rect 279451 65147 279499 65175
rect 279189 65113 279499 65147
rect 279189 65085 279237 65113
rect 279265 65085 279299 65113
rect 279327 65085 279361 65113
rect 279389 65085 279423 65113
rect 279451 65085 279499 65113
rect 279189 65051 279499 65085
rect 279189 65023 279237 65051
rect 279265 65023 279299 65051
rect 279327 65023 279361 65051
rect 279389 65023 279423 65051
rect 279451 65023 279499 65051
rect 279189 64989 279499 65023
rect 279189 64961 279237 64989
rect 279265 64961 279299 64989
rect 279327 64961 279361 64989
rect 279389 64961 279423 64989
rect 279451 64961 279499 64989
rect 276766 36577 276794 36582
rect 279189 56175 279499 64961
rect 279189 56147 279237 56175
rect 279265 56147 279299 56175
rect 279327 56147 279361 56175
rect 279389 56147 279423 56175
rect 279451 56147 279499 56175
rect 279189 56113 279499 56147
rect 279189 56085 279237 56113
rect 279265 56085 279299 56113
rect 279327 56085 279361 56113
rect 279389 56085 279423 56113
rect 279451 56085 279499 56113
rect 279189 56051 279499 56085
rect 279189 56023 279237 56051
rect 279265 56023 279299 56051
rect 279327 56023 279361 56051
rect 279389 56023 279423 56051
rect 279451 56023 279499 56051
rect 279189 55989 279499 56023
rect 279189 55961 279237 55989
rect 279265 55961 279299 55989
rect 279327 55961 279361 55989
rect 279389 55961 279423 55989
rect 279451 55961 279499 55989
rect 279189 47175 279499 55961
rect 279189 47147 279237 47175
rect 279265 47147 279299 47175
rect 279327 47147 279361 47175
rect 279389 47147 279423 47175
rect 279451 47147 279499 47175
rect 279189 47113 279499 47147
rect 279189 47085 279237 47113
rect 279265 47085 279299 47113
rect 279327 47085 279361 47113
rect 279389 47085 279423 47113
rect 279451 47085 279499 47113
rect 279189 47051 279499 47085
rect 279189 47023 279237 47051
rect 279265 47023 279299 47051
rect 279327 47023 279361 47051
rect 279389 47023 279423 47051
rect 279451 47023 279499 47051
rect 279189 46989 279499 47023
rect 279189 46961 279237 46989
rect 279265 46961 279299 46989
rect 279327 46961 279361 46989
rect 279389 46961 279423 46989
rect 279451 46961 279499 46989
rect 279189 38175 279499 46961
rect 279189 38147 279237 38175
rect 279265 38147 279299 38175
rect 279327 38147 279361 38175
rect 279389 38147 279423 38175
rect 279451 38147 279499 38175
rect 279189 38113 279499 38147
rect 279189 38085 279237 38113
rect 279265 38085 279299 38113
rect 279327 38085 279361 38113
rect 279389 38085 279423 38113
rect 279451 38085 279499 38113
rect 279189 38051 279499 38085
rect 279189 38023 279237 38051
rect 279265 38023 279299 38051
rect 279327 38023 279361 38051
rect 279389 38023 279423 38051
rect 279451 38023 279499 38051
rect 279189 37989 279499 38023
rect 279189 37961 279237 37989
rect 279265 37961 279299 37989
rect 279327 37961 279361 37989
rect 279389 37961 279423 37989
rect 279451 37961 279499 37989
rect 276094 23361 276122 23366
rect 279189 29175 279499 37961
rect 279189 29147 279237 29175
rect 279265 29147 279299 29175
rect 279327 29147 279361 29175
rect 279389 29147 279423 29175
rect 279451 29147 279499 29175
rect 279189 29113 279499 29147
rect 279189 29085 279237 29113
rect 279265 29085 279299 29113
rect 279327 29085 279361 29113
rect 279389 29085 279423 29113
rect 279451 29085 279499 29113
rect 279189 29051 279499 29085
rect 279189 29023 279237 29051
rect 279265 29023 279299 29051
rect 279327 29023 279361 29051
rect 279389 29023 279423 29051
rect 279451 29023 279499 29051
rect 279189 28989 279499 29023
rect 279189 28961 279237 28989
rect 279265 28961 279299 28989
rect 279327 28961 279361 28989
rect 279389 28961 279423 28989
rect 279451 28961 279499 28989
rect 275982 16809 276010 16814
rect 279189 20175 279499 28961
rect 279189 20147 279237 20175
rect 279265 20147 279299 20175
rect 279327 20147 279361 20175
rect 279389 20147 279423 20175
rect 279451 20147 279499 20175
rect 279189 20113 279499 20147
rect 279189 20085 279237 20113
rect 279265 20085 279299 20113
rect 279327 20085 279361 20113
rect 279389 20085 279423 20113
rect 279451 20085 279499 20113
rect 279189 20051 279499 20085
rect 279189 20023 279237 20051
rect 279265 20023 279299 20051
rect 279327 20023 279361 20051
rect 279389 20023 279423 20051
rect 279451 20023 279499 20051
rect 279189 19989 279499 20023
rect 279189 19961 279237 19989
rect 279265 19961 279299 19989
rect 279327 19961 279361 19989
rect 279389 19961 279423 19989
rect 279451 19961 279499 19989
rect 275926 3537 275954 3542
rect 279189 11175 279499 19961
rect 279189 11147 279237 11175
rect 279265 11147 279299 11175
rect 279327 11147 279361 11175
rect 279389 11147 279423 11175
rect 279451 11147 279499 11175
rect 279189 11113 279499 11147
rect 279189 11085 279237 11113
rect 279265 11085 279299 11113
rect 279327 11085 279361 11113
rect 279389 11085 279423 11113
rect 279451 11085 279499 11113
rect 279189 11051 279499 11085
rect 279189 11023 279237 11051
rect 279265 11023 279299 11051
rect 279327 11023 279361 11051
rect 279389 11023 279423 11051
rect 279451 11023 279499 11051
rect 279189 10989 279499 11023
rect 279189 10961 279237 10989
rect 279265 10961 279299 10989
rect 279327 10961 279361 10989
rect 279389 10961 279423 10989
rect 279451 10961 279499 10989
rect 265689 -588 265737 -560
rect 265765 -588 265799 -560
rect 265827 -588 265861 -560
rect 265889 -588 265923 -560
rect 265951 -588 265999 -560
rect 265689 -622 265999 -588
rect 265689 -650 265737 -622
rect 265765 -650 265799 -622
rect 265827 -650 265861 -622
rect 265889 -650 265923 -622
rect 265951 -650 265999 -622
rect 265689 -684 265999 -650
rect 265689 -712 265737 -684
rect 265765 -712 265799 -684
rect 265827 -712 265861 -684
rect 265889 -712 265923 -684
rect 265951 -712 265999 -684
rect 265689 -746 265999 -712
rect 265689 -774 265737 -746
rect 265765 -774 265799 -746
rect 265827 -774 265861 -746
rect 265889 -774 265923 -746
rect 265951 -774 265999 -746
rect 265689 -822 265999 -774
rect 279189 2175 279499 10961
rect 279189 2147 279237 2175
rect 279265 2147 279299 2175
rect 279327 2147 279361 2175
rect 279389 2147 279423 2175
rect 279451 2147 279499 2175
rect 279189 2113 279499 2147
rect 279189 2085 279237 2113
rect 279265 2085 279299 2113
rect 279327 2085 279361 2113
rect 279389 2085 279423 2113
rect 279451 2085 279499 2113
rect 279189 2051 279499 2085
rect 279189 2023 279237 2051
rect 279265 2023 279299 2051
rect 279327 2023 279361 2051
rect 279389 2023 279423 2051
rect 279451 2023 279499 2051
rect 279189 1989 279499 2023
rect 279189 1961 279237 1989
rect 279265 1961 279299 1989
rect 279327 1961 279361 1989
rect 279389 1961 279423 1989
rect 279451 1961 279499 1989
rect 279189 -80 279499 1961
rect 279189 -108 279237 -80
rect 279265 -108 279299 -80
rect 279327 -108 279361 -80
rect 279389 -108 279423 -80
rect 279451 -108 279499 -80
rect 279189 -142 279499 -108
rect 279189 -170 279237 -142
rect 279265 -170 279299 -142
rect 279327 -170 279361 -142
rect 279389 -170 279423 -142
rect 279451 -170 279499 -142
rect 279189 -204 279499 -170
rect 279189 -232 279237 -204
rect 279265 -232 279299 -204
rect 279327 -232 279361 -204
rect 279389 -232 279423 -204
rect 279451 -232 279499 -204
rect 279189 -266 279499 -232
rect 279189 -294 279237 -266
rect 279265 -294 279299 -266
rect 279327 -294 279361 -266
rect 279389 -294 279423 -266
rect 279451 -294 279499 -266
rect 279189 -822 279499 -294
rect 281049 299086 281359 299134
rect 281049 299058 281097 299086
rect 281125 299058 281159 299086
rect 281187 299058 281221 299086
rect 281249 299058 281283 299086
rect 281311 299058 281359 299086
rect 281049 299024 281359 299058
rect 281049 298996 281097 299024
rect 281125 298996 281159 299024
rect 281187 298996 281221 299024
rect 281249 298996 281283 299024
rect 281311 298996 281359 299024
rect 281049 298962 281359 298996
rect 281049 298934 281097 298962
rect 281125 298934 281159 298962
rect 281187 298934 281221 298962
rect 281249 298934 281283 298962
rect 281311 298934 281359 298962
rect 281049 298900 281359 298934
rect 281049 298872 281097 298900
rect 281125 298872 281159 298900
rect 281187 298872 281221 298900
rect 281249 298872 281283 298900
rect 281311 298872 281359 298900
rect 281049 293175 281359 298872
rect 281049 293147 281097 293175
rect 281125 293147 281159 293175
rect 281187 293147 281221 293175
rect 281249 293147 281283 293175
rect 281311 293147 281359 293175
rect 281049 293113 281359 293147
rect 281049 293085 281097 293113
rect 281125 293085 281159 293113
rect 281187 293085 281221 293113
rect 281249 293085 281283 293113
rect 281311 293085 281359 293113
rect 281049 293051 281359 293085
rect 281049 293023 281097 293051
rect 281125 293023 281159 293051
rect 281187 293023 281221 293051
rect 281249 293023 281283 293051
rect 281311 293023 281359 293051
rect 281049 292989 281359 293023
rect 281049 292961 281097 292989
rect 281125 292961 281159 292989
rect 281187 292961 281221 292989
rect 281249 292961 281283 292989
rect 281311 292961 281359 292989
rect 281049 284175 281359 292961
rect 281049 284147 281097 284175
rect 281125 284147 281159 284175
rect 281187 284147 281221 284175
rect 281249 284147 281283 284175
rect 281311 284147 281359 284175
rect 281049 284113 281359 284147
rect 281049 284085 281097 284113
rect 281125 284085 281159 284113
rect 281187 284085 281221 284113
rect 281249 284085 281283 284113
rect 281311 284085 281359 284113
rect 281049 284051 281359 284085
rect 281049 284023 281097 284051
rect 281125 284023 281159 284051
rect 281187 284023 281221 284051
rect 281249 284023 281283 284051
rect 281311 284023 281359 284051
rect 281049 283989 281359 284023
rect 281049 283961 281097 283989
rect 281125 283961 281159 283989
rect 281187 283961 281221 283989
rect 281249 283961 281283 283989
rect 281311 283961 281359 283989
rect 281049 275175 281359 283961
rect 281049 275147 281097 275175
rect 281125 275147 281159 275175
rect 281187 275147 281221 275175
rect 281249 275147 281283 275175
rect 281311 275147 281359 275175
rect 281049 275113 281359 275147
rect 281049 275085 281097 275113
rect 281125 275085 281159 275113
rect 281187 275085 281221 275113
rect 281249 275085 281283 275113
rect 281311 275085 281359 275113
rect 281049 275051 281359 275085
rect 281049 275023 281097 275051
rect 281125 275023 281159 275051
rect 281187 275023 281221 275051
rect 281249 275023 281283 275051
rect 281311 275023 281359 275051
rect 281049 274989 281359 275023
rect 281049 274961 281097 274989
rect 281125 274961 281159 274989
rect 281187 274961 281221 274989
rect 281249 274961 281283 274989
rect 281311 274961 281359 274989
rect 281049 266175 281359 274961
rect 281049 266147 281097 266175
rect 281125 266147 281159 266175
rect 281187 266147 281221 266175
rect 281249 266147 281283 266175
rect 281311 266147 281359 266175
rect 281049 266113 281359 266147
rect 281049 266085 281097 266113
rect 281125 266085 281159 266113
rect 281187 266085 281221 266113
rect 281249 266085 281283 266113
rect 281311 266085 281359 266113
rect 281049 266051 281359 266085
rect 281049 266023 281097 266051
rect 281125 266023 281159 266051
rect 281187 266023 281221 266051
rect 281249 266023 281283 266051
rect 281311 266023 281359 266051
rect 281049 265989 281359 266023
rect 281049 265961 281097 265989
rect 281125 265961 281159 265989
rect 281187 265961 281221 265989
rect 281249 265961 281283 265989
rect 281311 265961 281359 265989
rect 281049 257175 281359 265961
rect 281049 257147 281097 257175
rect 281125 257147 281159 257175
rect 281187 257147 281221 257175
rect 281249 257147 281283 257175
rect 281311 257147 281359 257175
rect 281049 257113 281359 257147
rect 281049 257085 281097 257113
rect 281125 257085 281159 257113
rect 281187 257085 281221 257113
rect 281249 257085 281283 257113
rect 281311 257085 281359 257113
rect 281049 257051 281359 257085
rect 281049 257023 281097 257051
rect 281125 257023 281159 257051
rect 281187 257023 281221 257051
rect 281249 257023 281283 257051
rect 281311 257023 281359 257051
rect 281049 256989 281359 257023
rect 281049 256961 281097 256989
rect 281125 256961 281159 256989
rect 281187 256961 281221 256989
rect 281249 256961 281283 256989
rect 281311 256961 281359 256989
rect 281049 248175 281359 256961
rect 281049 248147 281097 248175
rect 281125 248147 281159 248175
rect 281187 248147 281221 248175
rect 281249 248147 281283 248175
rect 281311 248147 281359 248175
rect 281049 248113 281359 248147
rect 281049 248085 281097 248113
rect 281125 248085 281159 248113
rect 281187 248085 281221 248113
rect 281249 248085 281283 248113
rect 281311 248085 281359 248113
rect 281049 248051 281359 248085
rect 281049 248023 281097 248051
rect 281125 248023 281159 248051
rect 281187 248023 281221 248051
rect 281249 248023 281283 248051
rect 281311 248023 281359 248051
rect 281049 247989 281359 248023
rect 281049 247961 281097 247989
rect 281125 247961 281159 247989
rect 281187 247961 281221 247989
rect 281249 247961 281283 247989
rect 281311 247961 281359 247989
rect 281049 239175 281359 247961
rect 281049 239147 281097 239175
rect 281125 239147 281159 239175
rect 281187 239147 281221 239175
rect 281249 239147 281283 239175
rect 281311 239147 281359 239175
rect 281049 239113 281359 239147
rect 281049 239085 281097 239113
rect 281125 239085 281159 239113
rect 281187 239085 281221 239113
rect 281249 239085 281283 239113
rect 281311 239085 281359 239113
rect 281049 239051 281359 239085
rect 281049 239023 281097 239051
rect 281125 239023 281159 239051
rect 281187 239023 281221 239051
rect 281249 239023 281283 239051
rect 281311 239023 281359 239051
rect 281049 238989 281359 239023
rect 281049 238961 281097 238989
rect 281125 238961 281159 238989
rect 281187 238961 281221 238989
rect 281249 238961 281283 238989
rect 281311 238961 281359 238989
rect 281049 230175 281359 238961
rect 281049 230147 281097 230175
rect 281125 230147 281159 230175
rect 281187 230147 281221 230175
rect 281249 230147 281283 230175
rect 281311 230147 281359 230175
rect 281049 230113 281359 230147
rect 281049 230085 281097 230113
rect 281125 230085 281159 230113
rect 281187 230085 281221 230113
rect 281249 230085 281283 230113
rect 281311 230085 281359 230113
rect 281049 230051 281359 230085
rect 281049 230023 281097 230051
rect 281125 230023 281159 230051
rect 281187 230023 281221 230051
rect 281249 230023 281283 230051
rect 281311 230023 281359 230051
rect 281049 229989 281359 230023
rect 281049 229961 281097 229989
rect 281125 229961 281159 229989
rect 281187 229961 281221 229989
rect 281249 229961 281283 229989
rect 281311 229961 281359 229989
rect 281049 221175 281359 229961
rect 281049 221147 281097 221175
rect 281125 221147 281159 221175
rect 281187 221147 281221 221175
rect 281249 221147 281283 221175
rect 281311 221147 281359 221175
rect 281049 221113 281359 221147
rect 281049 221085 281097 221113
rect 281125 221085 281159 221113
rect 281187 221085 281221 221113
rect 281249 221085 281283 221113
rect 281311 221085 281359 221113
rect 281049 221051 281359 221085
rect 281049 221023 281097 221051
rect 281125 221023 281159 221051
rect 281187 221023 281221 221051
rect 281249 221023 281283 221051
rect 281311 221023 281359 221051
rect 281049 220989 281359 221023
rect 281049 220961 281097 220989
rect 281125 220961 281159 220989
rect 281187 220961 281221 220989
rect 281249 220961 281283 220989
rect 281311 220961 281359 220989
rect 281049 212175 281359 220961
rect 281049 212147 281097 212175
rect 281125 212147 281159 212175
rect 281187 212147 281221 212175
rect 281249 212147 281283 212175
rect 281311 212147 281359 212175
rect 281049 212113 281359 212147
rect 281049 212085 281097 212113
rect 281125 212085 281159 212113
rect 281187 212085 281221 212113
rect 281249 212085 281283 212113
rect 281311 212085 281359 212113
rect 281049 212051 281359 212085
rect 281049 212023 281097 212051
rect 281125 212023 281159 212051
rect 281187 212023 281221 212051
rect 281249 212023 281283 212051
rect 281311 212023 281359 212051
rect 281049 211989 281359 212023
rect 281049 211961 281097 211989
rect 281125 211961 281159 211989
rect 281187 211961 281221 211989
rect 281249 211961 281283 211989
rect 281311 211961 281359 211989
rect 281049 203175 281359 211961
rect 281049 203147 281097 203175
rect 281125 203147 281159 203175
rect 281187 203147 281221 203175
rect 281249 203147 281283 203175
rect 281311 203147 281359 203175
rect 281049 203113 281359 203147
rect 281049 203085 281097 203113
rect 281125 203085 281159 203113
rect 281187 203085 281221 203113
rect 281249 203085 281283 203113
rect 281311 203085 281359 203113
rect 281049 203051 281359 203085
rect 281049 203023 281097 203051
rect 281125 203023 281159 203051
rect 281187 203023 281221 203051
rect 281249 203023 281283 203051
rect 281311 203023 281359 203051
rect 281049 202989 281359 203023
rect 281049 202961 281097 202989
rect 281125 202961 281159 202989
rect 281187 202961 281221 202989
rect 281249 202961 281283 202989
rect 281311 202961 281359 202989
rect 281049 194175 281359 202961
rect 281049 194147 281097 194175
rect 281125 194147 281159 194175
rect 281187 194147 281221 194175
rect 281249 194147 281283 194175
rect 281311 194147 281359 194175
rect 281049 194113 281359 194147
rect 281049 194085 281097 194113
rect 281125 194085 281159 194113
rect 281187 194085 281221 194113
rect 281249 194085 281283 194113
rect 281311 194085 281359 194113
rect 281049 194051 281359 194085
rect 281049 194023 281097 194051
rect 281125 194023 281159 194051
rect 281187 194023 281221 194051
rect 281249 194023 281283 194051
rect 281311 194023 281359 194051
rect 281049 193989 281359 194023
rect 281049 193961 281097 193989
rect 281125 193961 281159 193989
rect 281187 193961 281221 193989
rect 281249 193961 281283 193989
rect 281311 193961 281359 193989
rect 281049 185175 281359 193961
rect 281049 185147 281097 185175
rect 281125 185147 281159 185175
rect 281187 185147 281221 185175
rect 281249 185147 281283 185175
rect 281311 185147 281359 185175
rect 281049 185113 281359 185147
rect 281049 185085 281097 185113
rect 281125 185085 281159 185113
rect 281187 185085 281221 185113
rect 281249 185085 281283 185113
rect 281311 185085 281359 185113
rect 281049 185051 281359 185085
rect 281049 185023 281097 185051
rect 281125 185023 281159 185051
rect 281187 185023 281221 185051
rect 281249 185023 281283 185051
rect 281311 185023 281359 185051
rect 281049 184989 281359 185023
rect 281049 184961 281097 184989
rect 281125 184961 281159 184989
rect 281187 184961 281221 184989
rect 281249 184961 281283 184989
rect 281311 184961 281359 184989
rect 281049 176175 281359 184961
rect 281049 176147 281097 176175
rect 281125 176147 281159 176175
rect 281187 176147 281221 176175
rect 281249 176147 281283 176175
rect 281311 176147 281359 176175
rect 281049 176113 281359 176147
rect 281049 176085 281097 176113
rect 281125 176085 281159 176113
rect 281187 176085 281221 176113
rect 281249 176085 281283 176113
rect 281311 176085 281359 176113
rect 281049 176051 281359 176085
rect 281049 176023 281097 176051
rect 281125 176023 281159 176051
rect 281187 176023 281221 176051
rect 281249 176023 281283 176051
rect 281311 176023 281359 176051
rect 281049 175989 281359 176023
rect 281049 175961 281097 175989
rect 281125 175961 281159 175989
rect 281187 175961 281221 175989
rect 281249 175961 281283 175989
rect 281311 175961 281359 175989
rect 281049 167175 281359 175961
rect 281049 167147 281097 167175
rect 281125 167147 281159 167175
rect 281187 167147 281221 167175
rect 281249 167147 281283 167175
rect 281311 167147 281359 167175
rect 281049 167113 281359 167147
rect 281049 167085 281097 167113
rect 281125 167085 281159 167113
rect 281187 167085 281221 167113
rect 281249 167085 281283 167113
rect 281311 167085 281359 167113
rect 281049 167051 281359 167085
rect 281049 167023 281097 167051
rect 281125 167023 281159 167051
rect 281187 167023 281221 167051
rect 281249 167023 281283 167051
rect 281311 167023 281359 167051
rect 281049 166989 281359 167023
rect 281049 166961 281097 166989
rect 281125 166961 281159 166989
rect 281187 166961 281221 166989
rect 281249 166961 281283 166989
rect 281311 166961 281359 166989
rect 281049 158175 281359 166961
rect 281049 158147 281097 158175
rect 281125 158147 281159 158175
rect 281187 158147 281221 158175
rect 281249 158147 281283 158175
rect 281311 158147 281359 158175
rect 281049 158113 281359 158147
rect 281049 158085 281097 158113
rect 281125 158085 281159 158113
rect 281187 158085 281221 158113
rect 281249 158085 281283 158113
rect 281311 158085 281359 158113
rect 281049 158051 281359 158085
rect 281049 158023 281097 158051
rect 281125 158023 281159 158051
rect 281187 158023 281221 158051
rect 281249 158023 281283 158051
rect 281311 158023 281359 158051
rect 281049 157989 281359 158023
rect 281049 157961 281097 157989
rect 281125 157961 281159 157989
rect 281187 157961 281221 157989
rect 281249 157961 281283 157989
rect 281311 157961 281359 157989
rect 281049 149175 281359 157961
rect 281049 149147 281097 149175
rect 281125 149147 281159 149175
rect 281187 149147 281221 149175
rect 281249 149147 281283 149175
rect 281311 149147 281359 149175
rect 281049 149113 281359 149147
rect 281049 149085 281097 149113
rect 281125 149085 281159 149113
rect 281187 149085 281221 149113
rect 281249 149085 281283 149113
rect 281311 149085 281359 149113
rect 281049 149051 281359 149085
rect 281049 149023 281097 149051
rect 281125 149023 281159 149051
rect 281187 149023 281221 149051
rect 281249 149023 281283 149051
rect 281311 149023 281359 149051
rect 281049 148989 281359 149023
rect 281049 148961 281097 148989
rect 281125 148961 281159 148989
rect 281187 148961 281221 148989
rect 281249 148961 281283 148989
rect 281311 148961 281359 148989
rect 281049 140175 281359 148961
rect 281049 140147 281097 140175
rect 281125 140147 281159 140175
rect 281187 140147 281221 140175
rect 281249 140147 281283 140175
rect 281311 140147 281359 140175
rect 281049 140113 281359 140147
rect 281049 140085 281097 140113
rect 281125 140085 281159 140113
rect 281187 140085 281221 140113
rect 281249 140085 281283 140113
rect 281311 140085 281359 140113
rect 281049 140051 281359 140085
rect 281049 140023 281097 140051
rect 281125 140023 281159 140051
rect 281187 140023 281221 140051
rect 281249 140023 281283 140051
rect 281311 140023 281359 140051
rect 281049 139989 281359 140023
rect 281049 139961 281097 139989
rect 281125 139961 281159 139989
rect 281187 139961 281221 139989
rect 281249 139961 281283 139989
rect 281311 139961 281359 139989
rect 281049 131175 281359 139961
rect 281049 131147 281097 131175
rect 281125 131147 281159 131175
rect 281187 131147 281221 131175
rect 281249 131147 281283 131175
rect 281311 131147 281359 131175
rect 281049 131113 281359 131147
rect 281049 131085 281097 131113
rect 281125 131085 281159 131113
rect 281187 131085 281221 131113
rect 281249 131085 281283 131113
rect 281311 131085 281359 131113
rect 281049 131051 281359 131085
rect 281049 131023 281097 131051
rect 281125 131023 281159 131051
rect 281187 131023 281221 131051
rect 281249 131023 281283 131051
rect 281311 131023 281359 131051
rect 281049 130989 281359 131023
rect 281049 130961 281097 130989
rect 281125 130961 281159 130989
rect 281187 130961 281221 130989
rect 281249 130961 281283 130989
rect 281311 130961 281359 130989
rect 281049 122175 281359 130961
rect 281049 122147 281097 122175
rect 281125 122147 281159 122175
rect 281187 122147 281221 122175
rect 281249 122147 281283 122175
rect 281311 122147 281359 122175
rect 281049 122113 281359 122147
rect 281049 122085 281097 122113
rect 281125 122085 281159 122113
rect 281187 122085 281221 122113
rect 281249 122085 281283 122113
rect 281311 122085 281359 122113
rect 281049 122051 281359 122085
rect 281049 122023 281097 122051
rect 281125 122023 281159 122051
rect 281187 122023 281221 122051
rect 281249 122023 281283 122051
rect 281311 122023 281359 122051
rect 281049 121989 281359 122023
rect 281049 121961 281097 121989
rect 281125 121961 281159 121989
rect 281187 121961 281221 121989
rect 281249 121961 281283 121989
rect 281311 121961 281359 121989
rect 281049 113175 281359 121961
rect 281049 113147 281097 113175
rect 281125 113147 281159 113175
rect 281187 113147 281221 113175
rect 281249 113147 281283 113175
rect 281311 113147 281359 113175
rect 281049 113113 281359 113147
rect 281049 113085 281097 113113
rect 281125 113085 281159 113113
rect 281187 113085 281221 113113
rect 281249 113085 281283 113113
rect 281311 113085 281359 113113
rect 281049 113051 281359 113085
rect 281049 113023 281097 113051
rect 281125 113023 281159 113051
rect 281187 113023 281221 113051
rect 281249 113023 281283 113051
rect 281311 113023 281359 113051
rect 281049 112989 281359 113023
rect 281049 112961 281097 112989
rect 281125 112961 281159 112989
rect 281187 112961 281221 112989
rect 281249 112961 281283 112989
rect 281311 112961 281359 112989
rect 281049 104175 281359 112961
rect 281049 104147 281097 104175
rect 281125 104147 281159 104175
rect 281187 104147 281221 104175
rect 281249 104147 281283 104175
rect 281311 104147 281359 104175
rect 281049 104113 281359 104147
rect 281049 104085 281097 104113
rect 281125 104085 281159 104113
rect 281187 104085 281221 104113
rect 281249 104085 281283 104113
rect 281311 104085 281359 104113
rect 281049 104051 281359 104085
rect 281049 104023 281097 104051
rect 281125 104023 281159 104051
rect 281187 104023 281221 104051
rect 281249 104023 281283 104051
rect 281311 104023 281359 104051
rect 281049 103989 281359 104023
rect 281049 103961 281097 103989
rect 281125 103961 281159 103989
rect 281187 103961 281221 103989
rect 281249 103961 281283 103989
rect 281311 103961 281359 103989
rect 281049 95175 281359 103961
rect 281049 95147 281097 95175
rect 281125 95147 281159 95175
rect 281187 95147 281221 95175
rect 281249 95147 281283 95175
rect 281311 95147 281359 95175
rect 281049 95113 281359 95147
rect 281049 95085 281097 95113
rect 281125 95085 281159 95113
rect 281187 95085 281221 95113
rect 281249 95085 281283 95113
rect 281311 95085 281359 95113
rect 281049 95051 281359 95085
rect 281049 95023 281097 95051
rect 281125 95023 281159 95051
rect 281187 95023 281221 95051
rect 281249 95023 281283 95051
rect 281311 95023 281359 95051
rect 281049 94989 281359 95023
rect 281049 94961 281097 94989
rect 281125 94961 281159 94989
rect 281187 94961 281221 94989
rect 281249 94961 281283 94989
rect 281311 94961 281359 94989
rect 281049 86175 281359 94961
rect 281049 86147 281097 86175
rect 281125 86147 281159 86175
rect 281187 86147 281221 86175
rect 281249 86147 281283 86175
rect 281311 86147 281359 86175
rect 281049 86113 281359 86147
rect 281049 86085 281097 86113
rect 281125 86085 281159 86113
rect 281187 86085 281221 86113
rect 281249 86085 281283 86113
rect 281311 86085 281359 86113
rect 281049 86051 281359 86085
rect 281049 86023 281097 86051
rect 281125 86023 281159 86051
rect 281187 86023 281221 86051
rect 281249 86023 281283 86051
rect 281311 86023 281359 86051
rect 281049 85989 281359 86023
rect 281049 85961 281097 85989
rect 281125 85961 281159 85989
rect 281187 85961 281221 85989
rect 281249 85961 281283 85989
rect 281311 85961 281359 85989
rect 281049 77175 281359 85961
rect 281049 77147 281097 77175
rect 281125 77147 281159 77175
rect 281187 77147 281221 77175
rect 281249 77147 281283 77175
rect 281311 77147 281359 77175
rect 281049 77113 281359 77147
rect 281049 77085 281097 77113
rect 281125 77085 281159 77113
rect 281187 77085 281221 77113
rect 281249 77085 281283 77113
rect 281311 77085 281359 77113
rect 281049 77051 281359 77085
rect 281049 77023 281097 77051
rect 281125 77023 281159 77051
rect 281187 77023 281221 77051
rect 281249 77023 281283 77051
rect 281311 77023 281359 77051
rect 281049 76989 281359 77023
rect 281049 76961 281097 76989
rect 281125 76961 281159 76989
rect 281187 76961 281221 76989
rect 281249 76961 281283 76989
rect 281311 76961 281359 76989
rect 281049 68175 281359 76961
rect 281049 68147 281097 68175
rect 281125 68147 281159 68175
rect 281187 68147 281221 68175
rect 281249 68147 281283 68175
rect 281311 68147 281359 68175
rect 281049 68113 281359 68147
rect 281049 68085 281097 68113
rect 281125 68085 281159 68113
rect 281187 68085 281221 68113
rect 281249 68085 281283 68113
rect 281311 68085 281359 68113
rect 281049 68051 281359 68085
rect 281049 68023 281097 68051
rect 281125 68023 281159 68051
rect 281187 68023 281221 68051
rect 281249 68023 281283 68051
rect 281311 68023 281359 68051
rect 281049 67989 281359 68023
rect 281049 67961 281097 67989
rect 281125 67961 281159 67989
rect 281187 67961 281221 67989
rect 281249 67961 281283 67989
rect 281311 67961 281359 67989
rect 281049 59175 281359 67961
rect 281049 59147 281097 59175
rect 281125 59147 281159 59175
rect 281187 59147 281221 59175
rect 281249 59147 281283 59175
rect 281311 59147 281359 59175
rect 281049 59113 281359 59147
rect 281049 59085 281097 59113
rect 281125 59085 281159 59113
rect 281187 59085 281221 59113
rect 281249 59085 281283 59113
rect 281311 59085 281359 59113
rect 281049 59051 281359 59085
rect 281049 59023 281097 59051
rect 281125 59023 281159 59051
rect 281187 59023 281221 59051
rect 281249 59023 281283 59051
rect 281311 59023 281359 59051
rect 281049 58989 281359 59023
rect 281049 58961 281097 58989
rect 281125 58961 281159 58989
rect 281187 58961 281221 58989
rect 281249 58961 281283 58989
rect 281311 58961 281359 58989
rect 281049 50175 281359 58961
rect 281049 50147 281097 50175
rect 281125 50147 281159 50175
rect 281187 50147 281221 50175
rect 281249 50147 281283 50175
rect 281311 50147 281359 50175
rect 281049 50113 281359 50147
rect 281049 50085 281097 50113
rect 281125 50085 281159 50113
rect 281187 50085 281221 50113
rect 281249 50085 281283 50113
rect 281311 50085 281359 50113
rect 281049 50051 281359 50085
rect 281049 50023 281097 50051
rect 281125 50023 281159 50051
rect 281187 50023 281221 50051
rect 281249 50023 281283 50051
rect 281311 50023 281359 50051
rect 281049 49989 281359 50023
rect 281049 49961 281097 49989
rect 281125 49961 281159 49989
rect 281187 49961 281221 49989
rect 281249 49961 281283 49989
rect 281311 49961 281359 49989
rect 281049 41175 281359 49961
rect 281049 41147 281097 41175
rect 281125 41147 281159 41175
rect 281187 41147 281221 41175
rect 281249 41147 281283 41175
rect 281311 41147 281359 41175
rect 281049 41113 281359 41147
rect 281049 41085 281097 41113
rect 281125 41085 281159 41113
rect 281187 41085 281221 41113
rect 281249 41085 281283 41113
rect 281311 41085 281359 41113
rect 281049 41051 281359 41085
rect 281049 41023 281097 41051
rect 281125 41023 281159 41051
rect 281187 41023 281221 41051
rect 281249 41023 281283 41051
rect 281311 41023 281359 41051
rect 281049 40989 281359 41023
rect 281049 40961 281097 40989
rect 281125 40961 281159 40989
rect 281187 40961 281221 40989
rect 281249 40961 281283 40989
rect 281311 40961 281359 40989
rect 281049 32175 281359 40961
rect 281049 32147 281097 32175
rect 281125 32147 281159 32175
rect 281187 32147 281221 32175
rect 281249 32147 281283 32175
rect 281311 32147 281359 32175
rect 281049 32113 281359 32147
rect 281049 32085 281097 32113
rect 281125 32085 281159 32113
rect 281187 32085 281221 32113
rect 281249 32085 281283 32113
rect 281311 32085 281359 32113
rect 281049 32051 281359 32085
rect 281049 32023 281097 32051
rect 281125 32023 281159 32051
rect 281187 32023 281221 32051
rect 281249 32023 281283 32051
rect 281311 32023 281359 32051
rect 281049 31989 281359 32023
rect 281049 31961 281097 31989
rect 281125 31961 281159 31989
rect 281187 31961 281221 31989
rect 281249 31961 281283 31989
rect 281311 31961 281359 31989
rect 281049 23175 281359 31961
rect 281049 23147 281097 23175
rect 281125 23147 281159 23175
rect 281187 23147 281221 23175
rect 281249 23147 281283 23175
rect 281311 23147 281359 23175
rect 281049 23113 281359 23147
rect 281049 23085 281097 23113
rect 281125 23085 281159 23113
rect 281187 23085 281221 23113
rect 281249 23085 281283 23113
rect 281311 23085 281359 23113
rect 281049 23051 281359 23085
rect 281049 23023 281097 23051
rect 281125 23023 281159 23051
rect 281187 23023 281221 23051
rect 281249 23023 281283 23051
rect 281311 23023 281359 23051
rect 281049 22989 281359 23023
rect 281049 22961 281097 22989
rect 281125 22961 281159 22989
rect 281187 22961 281221 22989
rect 281249 22961 281283 22989
rect 281311 22961 281359 22989
rect 281049 14175 281359 22961
rect 281049 14147 281097 14175
rect 281125 14147 281159 14175
rect 281187 14147 281221 14175
rect 281249 14147 281283 14175
rect 281311 14147 281359 14175
rect 281049 14113 281359 14147
rect 281049 14085 281097 14113
rect 281125 14085 281159 14113
rect 281187 14085 281221 14113
rect 281249 14085 281283 14113
rect 281311 14085 281359 14113
rect 281049 14051 281359 14085
rect 281049 14023 281097 14051
rect 281125 14023 281159 14051
rect 281187 14023 281221 14051
rect 281249 14023 281283 14051
rect 281311 14023 281359 14051
rect 281049 13989 281359 14023
rect 281049 13961 281097 13989
rect 281125 13961 281159 13989
rect 281187 13961 281221 13989
rect 281249 13961 281283 13989
rect 281311 13961 281359 13989
rect 281049 5175 281359 13961
rect 281049 5147 281097 5175
rect 281125 5147 281159 5175
rect 281187 5147 281221 5175
rect 281249 5147 281283 5175
rect 281311 5147 281359 5175
rect 281049 5113 281359 5147
rect 281049 5085 281097 5113
rect 281125 5085 281159 5113
rect 281187 5085 281221 5113
rect 281249 5085 281283 5113
rect 281311 5085 281359 5113
rect 281049 5051 281359 5085
rect 281049 5023 281097 5051
rect 281125 5023 281159 5051
rect 281187 5023 281221 5051
rect 281249 5023 281283 5051
rect 281311 5023 281359 5051
rect 281049 4989 281359 5023
rect 281049 4961 281097 4989
rect 281125 4961 281159 4989
rect 281187 4961 281221 4989
rect 281249 4961 281283 4989
rect 281311 4961 281359 4989
rect 281049 -560 281359 4961
rect 281049 -588 281097 -560
rect 281125 -588 281159 -560
rect 281187 -588 281221 -560
rect 281249 -588 281283 -560
rect 281311 -588 281359 -560
rect 281049 -622 281359 -588
rect 281049 -650 281097 -622
rect 281125 -650 281159 -622
rect 281187 -650 281221 -622
rect 281249 -650 281283 -622
rect 281311 -650 281359 -622
rect 281049 -684 281359 -650
rect 281049 -712 281097 -684
rect 281125 -712 281159 -684
rect 281187 -712 281221 -684
rect 281249 -712 281283 -684
rect 281311 -712 281359 -684
rect 281049 -746 281359 -712
rect 281049 -774 281097 -746
rect 281125 -774 281159 -746
rect 281187 -774 281221 -746
rect 281249 -774 281283 -746
rect 281311 -774 281359 -746
rect 281049 -822 281359 -774
rect 294549 298606 294859 299134
rect 294549 298578 294597 298606
rect 294625 298578 294659 298606
rect 294687 298578 294721 298606
rect 294749 298578 294783 298606
rect 294811 298578 294859 298606
rect 294549 298544 294859 298578
rect 294549 298516 294597 298544
rect 294625 298516 294659 298544
rect 294687 298516 294721 298544
rect 294749 298516 294783 298544
rect 294811 298516 294859 298544
rect 294549 298482 294859 298516
rect 294549 298454 294597 298482
rect 294625 298454 294659 298482
rect 294687 298454 294721 298482
rect 294749 298454 294783 298482
rect 294811 298454 294859 298482
rect 294549 298420 294859 298454
rect 294549 298392 294597 298420
rect 294625 298392 294659 298420
rect 294687 298392 294721 298420
rect 294749 298392 294783 298420
rect 294811 298392 294859 298420
rect 294549 290175 294859 298392
rect 294549 290147 294597 290175
rect 294625 290147 294659 290175
rect 294687 290147 294721 290175
rect 294749 290147 294783 290175
rect 294811 290147 294859 290175
rect 294549 290113 294859 290147
rect 294549 290085 294597 290113
rect 294625 290085 294659 290113
rect 294687 290085 294721 290113
rect 294749 290085 294783 290113
rect 294811 290085 294859 290113
rect 294549 290051 294859 290085
rect 294549 290023 294597 290051
rect 294625 290023 294659 290051
rect 294687 290023 294721 290051
rect 294749 290023 294783 290051
rect 294811 290023 294859 290051
rect 294549 289989 294859 290023
rect 294549 289961 294597 289989
rect 294625 289961 294659 289989
rect 294687 289961 294721 289989
rect 294749 289961 294783 289989
rect 294811 289961 294859 289989
rect 294549 281175 294859 289961
rect 294549 281147 294597 281175
rect 294625 281147 294659 281175
rect 294687 281147 294721 281175
rect 294749 281147 294783 281175
rect 294811 281147 294859 281175
rect 294549 281113 294859 281147
rect 294549 281085 294597 281113
rect 294625 281085 294659 281113
rect 294687 281085 294721 281113
rect 294749 281085 294783 281113
rect 294811 281085 294859 281113
rect 296409 299086 296719 299134
rect 296409 299058 296457 299086
rect 296485 299058 296519 299086
rect 296547 299058 296581 299086
rect 296609 299058 296643 299086
rect 296671 299058 296719 299086
rect 296409 299024 296719 299058
rect 296409 298996 296457 299024
rect 296485 298996 296519 299024
rect 296547 298996 296581 299024
rect 296609 298996 296643 299024
rect 296671 298996 296719 299024
rect 296409 298962 296719 298996
rect 296409 298934 296457 298962
rect 296485 298934 296519 298962
rect 296547 298934 296581 298962
rect 296609 298934 296643 298962
rect 296671 298934 296719 298962
rect 296409 298900 296719 298934
rect 296409 298872 296457 298900
rect 296485 298872 296519 298900
rect 296547 298872 296581 298900
rect 296609 298872 296643 298900
rect 296671 298872 296719 298900
rect 296409 293175 296719 298872
rect 298680 299086 298990 299134
rect 298680 299058 298728 299086
rect 298756 299058 298790 299086
rect 298818 299058 298852 299086
rect 298880 299058 298914 299086
rect 298942 299058 298990 299086
rect 298680 299024 298990 299058
rect 298680 298996 298728 299024
rect 298756 298996 298790 299024
rect 298818 298996 298852 299024
rect 298880 298996 298914 299024
rect 298942 298996 298990 299024
rect 298680 298962 298990 298996
rect 298680 298934 298728 298962
rect 298756 298934 298790 298962
rect 298818 298934 298852 298962
rect 298880 298934 298914 298962
rect 298942 298934 298990 298962
rect 298680 298900 298990 298934
rect 298680 298872 298728 298900
rect 298756 298872 298790 298900
rect 298818 298872 298852 298900
rect 298880 298872 298914 298900
rect 298942 298872 298990 298900
rect 296409 293147 296457 293175
rect 296485 293147 296519 293175
rect 296547 293147 296581 293175
rect 296609 293147 296643 293175
rect 296671 293147 296719 293175
rect 296409 293113 296719 293147
rect 296409 293085 296457 293113
rect 296485 293085 296519 293113
rect 296547 293085 296581 293113
rect 296609 293085 296643 293113
rect 296671 293085 296719 293113
rect 296409 293051 296719 293085
rect 296409 293023 296457 293051
rect 296485 293023 296519 293051
rect 296547 293023 296581 293051
rect 296609 293023 296643 293051
rect 296671 293023 296719 293051
rect 296409 292989 296719 293023
rect 296409 292961 296457 292989
rect 296485 292961 296519 292989
rect 296547 292961 296581 292989
rect 296609 292961 296643 292989
rect 296671 292961 296719 292989
rect 296409 284175 296719 292961
rect 296409 284147 296457 284175
rect 296485 284147 296519 284175
rect 296547 284147 296581 284175
rect 296609 284147 296643 284175
rect 296671 284147 296719 284175
rect 296409 284113 296719 284147
rect 296409 284085 296457 284113
rect 296485 284085 296519 284113
rect 296547 284085 296581 284113
rect 296609 284085 296643 284113
rect 296671 284085 296719 284113
rect 296409 284051 296719 284085
rect 296409 284023 296457 284051
rect 296485 284023 296519 284051
rect 296547 284023 296581 284051
rect 296609 284023 296643 284051
rect 296671 284023 296719 284051
rect 296409 283989 296719 284023
rect 296409 283961 296457 283989
rect 296485 283961 296519 283989
rect 296547 283961 296581 283989
rect 296609 283961 296643 283989
rect 296671 283961 296719 283989
rect 294549 281051 294859 281085
rect 294549 281023 294597 281051
rect 294625 281023 294659 281051
rect 294687 281023 294721 281051
rect 294749 281023 294783 281051
rect 294811 281023 294859 281051
rect 294549 280989 294859 281023
rect 294549 280961 294597 280989
rect 294625 280961 294659 280989
rect 294687 280961 294721 280989
rect 294749 280961 294783 280989
rect 294811 280961 294859 280989
rect 294549 272175 294859 280961
rect 294549 272147 294597 272175
rect 294625 272147 294659 272175
rect 294687 272147 294721 272175
rect 294749 272147 294783 272175
rect 294811 272147 294859 272175
rect 294549 272113 294859 272147
rect 294549 272085 294597 272113
rect 294625 272085 294659 272113
rect 294687 272085 294721 272113
rect 294749 272085 294783 272113
rect 294811 272085 294859 272113
rect 294549 272051 294859 272085
rect 294549 272023 294597 272051
rect 294625 272023 294659 272051
rect 294687 272023 294721 272051
rect 294749 272023 294783 272051
rect 294811 272023 294859 272051
rect 294549 271989 294859 272023
rect 294549 271961 294597 271989
rect 294625 271961 294659 271989
rect 294687 271961 294721 271989
rect 294749 271961 294783 271989
rect 294811 271961 294859 271989
rect 294549 263175 294859 271961
rect 294549 263147 294597 263175
rect 294625 263147 294659 263175
rect 294687 263147 294721 263175
rect 294749 263147 294783 263175
rect 294811 263147 294859 263175
rect 294549 263113 294859 263147
rect 294549 263085 294597 263113
rect 294625 263085 294659 263113
rect 294687 263085 294721 263113
rect 294749 263085 294783 263113
rect 294811 263085 294859 263113
rect 294549 263051 294859 263085
rect 294549 263023 294597 263051
rect 294625 263023 294659 263051
rect 294687 263023 294721 263051
rect 294749 263023 294783 263051
rect 294811 263023 294859 263051
rect 294549 262989 294859 263023
rect 294549 262961 294597 262989
rect 294625 262961 294659 262989
rect 294687 262961 294721 262989
rect 294749 262961 294783 262989
rect 294811 262961 294859 262989
rect 294549 254175 294859 262961
rect 294549 254147 294597 254175
rect 294625 254147 294659 254175
rect 294687 254147 294721 254175
rect 294749 254147 294783 254175
rect 294811 254147 294859 254175
rect 294549 254113 294859 254147
rect 294549 254085 294597 254113
rect 294625 254085 294659 254113
rect 294687 254085 294721 254113
rect 294749 254085 294783 254113
rect 294811 254085 294859 254113
rect 294549 254051 294859 254085
rect 294549 254023 294597 254051
rect 294625 254023 294659 254051
rect 294687 254023 294721 254051
rect 294749 254023 294783 254051
rect 294811 254023 294859 254051
rect 294549 253989 294859 254023
rect 294549 253961 294597 253989
rect 294625 253961 294659 253989
rect 294687 253961 294721 253989
rect 294749 253961 294783 253989
rect 294811 253961 294859 253989
rect 294549 245175 294859 253961
rect 294549 245147 294597 245175
rect 294625 245147 294659 245175
rect 294687 245147 294721 245175
rect 294749 245147 294783 245175
rect 294811 245147 294859 245175
rect 294549 245113 294859 245147
rect 294549 245085 294597 245113
rect 294625 245085 294659 245113
rect 294687 245085 294721 245113
rect 294749 245085 294783 245113
rect 294811 245085 294859 245113
rect 294549 245051 294859 245085
rect 294549 245023 294597 245051
rect 294625 245023 294659 245051
rect 294687 245023 294721 245051
rect 294749 245023 294783 245051
rect 294811 245023 294859 245051
rect 294549 244989 294859 245023
rect 294549 244961 294597 244989
rect 294625 244961 294659 244989
rect 294687 244961 294721 244989
rect 294749 244961 294783 244989
rect 294811 244961 294859 244989
rect 294549 236175 294859 244961
rect 294549 236147 294597 236175
rect 294625 236147 294659 236175
rect 294687 236147 294721 236175
rect 294749 236147 294783 236175
rect 294811 236147 294859 236175
rect 294549 236113 294859 236147
rect 294549 236085 294597 236113
rect 294625 236085 294659 236113
rect 294687 236085 294721 236113
rect 294749 236085 294783 236113
rect 294811 236085 294859 236113
rect 294549 236051 294859 236085
rect 294549 236023 294597 236051
rect 294625 236023 294659 236051
rect 294687 236023 294721 236051
rect 294749 236023 294783 236051
rect 294811 236023 294859 236051
rect 294549 235989 294859 236023
rect 294549 235961 294597 235989
rect 294625 235961 294659 235989
rect 294687 235961 294721 235989
rect 294749 235961 294783 235989
rect 294811 235961 294859 235989
rect 294549 227175 294859 235961
rect 294549 227147 294597 227175
rect 294625 227147 294659 227175
rect 294687 227147 294721 227175
rect 294749 227147 294783 227175
rect 294811 227147 294859 227175
rect 294549 227113 294859 227147
rect 294549 227085 294597 227113
rect 294625 227085 294659 227113
rect 294687 227085 294721 227113
rect 294749 227085 294783 227113
rect 294811 227085 294859 227113
rect 294549 227051 294859 227085
rect 294549 227023 294597 227051
rect 294625 227023 294659 227051
rect 294687 227023 294721 227051
rect 294749 227023 294783 227051
rect 294811 227023 294859 227051
rect 294549 226989 294859 227023
rect 294549 226961 294597 226989
rect 294625 226961 294659 226989
rect 294687 226961 294721 226989
rect 294749 226961 294783 226989
rect 294811 226961 294859 226989
rect 294549 218175 294859 226961
rect 294549 218147 294597 218175
rect 294625 218147 294659 218175
rect 294687 218147 294721 218175
rect 294749 218147 294783 218175
rect 294811 218147 294859 218175
rect 294549 218113 294859 218147
rect 294549 218085 294597 218113
rect 294625 218085 294659 218113
rect 294687 218085 294721 218113
rect 294749 218085 294783 218113
rect 294811 218085 294859 218113
rect 294549 218051 294859 218085
rect 294549 218023 294597 218051
rect 294625 218023 294659 218051
rect 294687 218023 294721 218051
rect 294749 218023 294783 218051
rect 294811 218023 294859 218051
rect 294549 217989 294859 218023
rect 294549 217961 294597 217989
rect 294625 217961 294659 217989
rect 294687 217961 294721 217989
rect 294749 217961 294783 217989
rect 294811 217961 294859 217989
rect 294549 209175 294859 217961
rect 294549 209147 294597 209175
rect 294625 209147 294659 209175
rect 294687 209147 294721 209175
rect 294749 209147 294783 209175
rect 294811 209147 294859 209175
rect 294549 209113 294859 209147
rect 294549 209085 294597 209113
rect 294625 209085 294659 209113
rect 294687 209085 294721 209113
rect 294749 209085 294783 209113
rect 294811 209085 294859 209113
rect 294549 209051 294859 209085
rect 294549 209023 294597 209051
rect 294625 209023 294659 209051
rect 294687 209023 294721 209051
rect 294749 209023 294783 209051
rect 294811 209023 294859 209051
rect 294549 208989 294859 209023
rect 294549 208961 294597 208989
rect 294625 208961 294659 208989
rect 294687 208961 294721 208989
rect 294749 208961 294783 208989
rect 294811 208961 294859 208989
rect 294549 200175 294859 208961
rect 294549 200147 294597 200175
rect 294625 200147 294659 200175
rect 294687 200147 294721 200175
rect 294749 200147 294783 200175
rect 294811 200147 294859 200175
rect 294549 200113 294859 200147
rect 294549 200085 294597 200113
rect 294625 200085 294659 200113
rect 294687 200085 294721 200113
rect 294749 200085 294783 200113
rect 294811 200085 294859 200113
rect 294549 200051 294859 200085
rect 294549 200023 294597 200051
rect 294625 200023 294659 200051
rect 294687 200023 294721 200051
rect 294749 200023 294783 200051
rect 294811 200023 294859 200051
rect 294549 199989 294859 200023
rect 294549 199961 294597 199989
rect 294625 199961 294659 199989
rect 294687 199961 294721 199989
rect 294749 199961 294783 199989
rect 294811 199961 294859 199989
rect 294549 191175 294859 199961
rect 294549 191147 294597 191175
rect 294625 191147 294659 191175
rect 294687 191147 294721 191175
rect 294749 191147 294783 191175
rect 294811 191147 294859 191175
rect 294549 191113 294859 191147
rect 294549 191085 294597 191113
rect 294625 191085 294659 191113
rect 294687 191085 294721 191113
rect 294749 191085 294783 191113
rect 294811 191085 294859 191113
rect 294549 191051 294859 191085
rect 294549 191023 294597 191051
rect 294625 191023 294659 191051
rect 294687 191023 294721 191051
rect 294749 191023 294783 191051
rect 294811 191023 294859 191051
rect 294549 190989 294859 191023
rect 294549 190961 294597 190989
rect 294625 190961 294659 190989
rect 294687 190961 294721 190989
rect 294749 190961 294783 190989
rect 294811 190961 294859 190989
rect 294549 182175 294859 190961
rect 294549 182147 294597 182175
rect 294625 182147 294659 182175
rect 294687 182147 294721 182175
rect 294749 182147 294783 182175
rect 294811 182147 294859 182175
rect 294549 182113 294859 182147
rect 294549 182085 294597 182113
rect 294625 182085 294659 182113
rect 294687 182085 294721 182113
rect 294749 182085 294783 182113
rect 294811 182085 294859 182113
rect 294549 182051 294859 182085
rect 294549 182023 294597 182051
rect 294625 182023 294659 182051
rect 294687 182023 294721 182051
rect 294749 182023 294783 182051
rect 294811 182023 294859 182051
rect 294549 181989 294859 182023
rect 294549 181961 294597 181989
rect 294625 181961 294659 181989
rect 294687 181961 294721 181989
rect 294749 181961 294783 181989
rect 294811 181961 294859 181989
rect 294549 173175 294859 181961
rect 294549 173147 294597 173175
rect 294625 173147 294659 173175
rect 294687 173147 294721 173175
rect 294749 173147 294783 173175
rect 294811 173147 294859 173175
rect 294549 173113 294859 173147
rect 294549 173085 294597 173113
rect 294625 173085 294659 173113
rect 294687 173085 294721 173113
rect 294749 173085 294783 173113
rect 294811 173085 294859 173113
rect 294549 173051 294859 173085
rect 294549 173023 294597 173051
rect 294625 173023 294659 173051
rect 294687 173023 294721 173051
rect 294749 173023 294783 173051
rect 294811 173023 294859 173051
rect 294549 172989 294859 173023
rect 294549 172961 294597 172989
rect 294625 172961 294659 172989
rect 294687 172961 294721 172989
rect 294749 172961 294783 172989
rect 294811 172961 294859 172989
rect 294549 164175 294859 172961
rect 294549 164147 294597 164175
rect 294625 164147 294659 164175
rect 294687 164147 294721 164175
rect 294749 164147 294783 164175
rect 294811 164147 294859 164175
rect 294549 164113 294859 164147
rect 294549 164085 294597 164113
rect 294625 164085 294659 164113
rect 294687 164085 294721 164113
rect 294749 164085 294783 164113
rect 294811 164085 294859 164113
rect 294549 164051 294859 164085
rect 294549 164023 294597 164051
rect 294625 164023 294659 164051
rect 294687 164023 294721 164051
rect 294749 164023 294783 164051
rect 294811 164023 294859 164051
rect 294549 163989 294859 164023
rect 294549 163961 294597 163989
rect 294625 163961 294659 163989
rect 294687 163961 294721 163989
rect 294749 163961 294783 163989
rect 294811 163961 294859 163989
rect 294549 155175 294859 163961
rect 295246 281106 295274 281111
rect 295246 156786 295274 281078
rect 296409 275175 296719 283961
rect 296409 275147 296457 275175
rect 296485 275147 296519 275175
rect 296547 275147 296581 275175
rect 296609 275147 296643 275175
rect 296671 275147 296719 275175
rect 296409 275113 296719 275147
rect 296409 275085 296457 275113
rect 296485 275085 296519 275113
rect 296547 275085 296581 275113
rect 296609 275085 296643 275113
rect 296671 275085 296719 275113
rect 296409 275051 296719 275085
rect 296409 275023 296457 275051
rect 296485 275023 296519 275051
rect 296547 275023 296581 275051
rect 296609 275023 296643 275051
rect 296671 275023 296719 275051
rect 296409 274989 296719 275023
rect 296409 274961 296457 274989
rect 296485 274961 296519 274989
rect 296547 274961 296581 274989
rect 296609 274961 296643 274989
rect 296671 274961 296719 274989
rect 296409 266175 296719 274961
rect 296409 266147 296457 266175
rect 296485 266147 296519 266175
rect 296547 266147 296581 266175
rect 296609 266147 296643 266175
rect 296671 266147 296719 266175
rect 296409 266113 296719 266147
rect 296409 266085 296457 266113
rect 296485 266085 296519 266113
rect 296547 266085 296581 266113
rect 296609 266085 296643 266113
rect 296671 266085 296719 266113
rect 296409 266051 296719 266085
rect 296409 266023 296457 266051
rect 296485 266023 296519 266051
rect 296547 266023 296581 266051
rect 296609 266023 296643 266051
rect 296671 266023 296719 266051
rect 296409 265989 296719 266023
rect 296409 265961 296457 265989
rect 296485 265961 296519 265989
rect 296547 265961 296581 265989
rect 296609 265961 296643 265989
rect 296671 265961 296719 265989
rect 295246 156753 295274 156758
rect 295302 261282 295330 261287
rect 295302 155442 295330 261254
rect 296409 257175 296719 265961
rect 296409 257147 296457 257175
rect 296485 257147 296519 257175
rect 296547 257147 296581 257175
rect 296609 257147 296643 257175
rect 296671 257147 296719 257175
rect 296409 257113 296719 257147
rect 296409 257085 296457 257113
rect 296485 257085 296519 257113
rect 296547 257085 296581 257113
rect 296609 257085 296643 257113
rect 296671 257085 296719 257113
rect 296409 257051 296719 257085
rect 296409 257023 296457 257051
rect 296485 257023 296519 257051
rect 296547 257023 296581 257051
rect 296609 257023 296643 257051
rect 296671 257023 296719 257051
rect 296409 256989 296719 257023
rect 296409 256961 296457 256989
rect 296485 256961 296519 256989
rect 296547 256961 296581 256989
rect 296609 256961 296643 256989
rect 296671 256961 296719 256989
rect 296409 248175 296719 256961
rect 296409 248147 296457 248175
rect 296485 248147 296519 248175
rect 296547 248147 296581 248175
rect 296609 248147 296643 248175
rect 296671 248147 296719 248175
rect 296409 248113 296719 248147
rect 296409 248085 296457 248113
rect 296485 248085 296519 248113
rect 296547 248085 296581 248113
rect 296609 248085 296643 248113
rect 296671 248085 296719 248113
rect 296409 248051 296719 248085
rect 296409 248023 296457 248051
rect 296485 248023 296519 248051
rect 296547 248023 296581 248051
rect 296609 248023 296643 248051
rect 296671 248023 296719 248051
rect 296409 247989 296719 248023
rect 296409 247961 296457 247989
rect 296485 247961 296519 247989
rect 296547 247961 296581 247989
rect 296609 247961 296643 247989
rect 296671 247961 296719 247989
rect 295302 155409 295330 155414
rect 295358 241458 295386 241463
rect 294549 155147 294597 155175
rect 294625 155147 294659 155175
rect 294687 155147 294721 155175
rect 294749 155147 294783 155175
rect 294811 155147 294859 155175
rect 294549 155113 294859 155147
rect 294549 155085 294597 155113
rect 294625 155085 294659 155113
rect 294687 155085 294721 155113
rect 294749 155085 294783 155113
rect 294811 155085 294859 155113
rect 294549 155051 294859 155085
rect 294549 155023 294597 155051
rect 294625 155023 294659 155051
rect 294687 155023 294721 155051
rect 294749 155023 294783 155051
rect 294811 155023 294859 155051
rect 294549 154989 294859 155023
rect 294549 154961 294597 154989
rect 294625 154961 294659 154989
rect 294687 154961 294721 154989
rect 294749 154961 294783 154989
rect 294811 154961 294859 154989
rect 294549 146175 294859 154961
rect 295358 154098 295386 241430
rect 296409 239175 296719 247961
rect 296409 239147 296457 239175
rect 296485 239147 296519 239175
rect 296547 239147 296581 239175
rect 296609 239147 296643 239175
rect 296671 239147 296719 239175
rect 296409 239113 296719 239147
rect 296409 239085 296457 239113
rect 296485 239085 296519 239113
rect 296547 239085 296581 239113
rect 296609 239085 296643 239113
rect 296671 239085 296719 239113
rect 296409 239051 296719 239085
rect 296409 239023 296457 239051
rect 296485 239023 296519 239051
rect 296547 239023 296581 239051
rect 296609 239023 296643 239051
rect 296671 239023 296719 239051
rect 296409 238989 296719 239023
rect 296409 238961 296457 238989
rect 296485 238961 296519 238989
rect 296547 238961 296581 238989
rect 296609 238961 296643 238989
rect 296671 238961 296719 238989
rect 296409 230175 296719 238961
rect 296409 230147 296457 230175
rect 296485 230147 296519 230175
rect 296547 230147 296581 230175
rect 296609 230147 296643 230175
rect 296671 230147 296719 230175
rect 296409 230113 296719 230147
rect 296409 230085 296457 230113
rect 296485 230085 296519 230113
rect 296547 230085 296581 230113
rect 296609 230085 296643 230113
rect 296671 230085 296719 230113
rect 296409 230051 296719 230085
rect 296409 230023 296457 230051
rect 296485 230023 296519 230051
rect 296547 230023 296581 230051
rect 296609 230023 296643 230051
rect 296671 230023 296719 230051
rect 296409 229989 296719 230023
rect 296409 229961 296457 229989
rect 296485 229961 296519 229989
rect 296547 229961 296581 229989
rect 296609 229961 296643 229989
rect 296671 229961 296719 229989
rect 295358 154065 295386 154070
rect 295414 221634 295442 221639
rect 295414 152754 295442 221606
rect 296409 221175 296719 229961
rect 296409 221147 296457 221175
rect 296485 221147 296519 221175
rect 296547 221147 296581 221175
rect 296609 221147 296643 221175
rect 296671 221147 296719 221175
rect 296409 221113 296719 221147
rect 296409 221085 296457 221113
rect 296485 221085 296519 221113
rect 296547 221085 296581 221113
rect 296609 221085 296643 221113
rect 296671 221085 296719 221113
rect 296409 221051 296719 221085
rect 296409 221023 296457 221051
rect 296485 221023 296519 221051
rect 296547 221023 296581 221051
rect 296609 221023 296643 221051
rect 296671 221023 296719 221051
rect 296409 220989 296719 221023
rect 296409 220961 296457 220989
rect 296485 220961 296519 220989
rect 296547 220961 296581 220989
rect 296609 220961 296643 220989
rect 296671 220961 296719 220989
rect 296409 212175 296719 220961
rect 296409 212147 296457 212175
rect 296485 212147 296519 212175
rect 296547 212147 296581 212175
rect 296609 212147 296643 212175
rect 296671 212147 296719 212175
rect 296409 212113 296719 212147
rect 296409 212085 296457 212113
rect 296485 212085 296519 212113
rect 296547 212085 296581 212113
rect 296609 212085 296643 212113
rect 296671 212085 296719 212113
rect 296409 212051 296719 212085
rect 296409 212023 296457 212051
rect 296485 212023 296519 212051
rect 296547 212023 296581 212051
rect 296609 212023 296643 212051
rect 296671 212023 296719 212051
rect 296409 211989 296719 212023
rect 296409 211961 296457 211989
rect 296485 211961 296519 211989
rect 296547 211961 296581 211989
rect 296609 211961 296643 211989
rect 296671 211961 296719 211989
rect 296409 203175 296719 211961
rect 296409 203147 296457 203175
rect 296485 203147 296519 203175
rect 296547 203147 296581 203175
rect 296609 203147 296643 203175
rect 296671 203147 296719 203175
rect 296409 203113 296719 203147
rect 296409 203085 296457 203113
rect 296485 203085 296519 203113
rect 296547 203085 296581 203113
rect 296609 203085 296643 203113
rect 296671 203085 296719 203113
rect 296409 203051 296719 203085
rect 296409 203023 296457 203051
rect 296485 203023 296519 203051
rect 296547 203023 296581 203051
rect 296609 203023 296643 203051
rect 296671 203023 296719 203051
rect 296409 202989 296719 203023
rect 296409 202961 296457 202989
rect 296485 202961 296519 202989
rect 296547 202961 296581 202989
rect 296609 202961 296643 202989
rect 296671 202961 296719 202989
rect 295414 152721 295442 152726
rect 295470 201810 295498 201815
rect 295470 151410 295498 201782
rect 295470 151377 295498 151382
rect 296409 194175 296719 202961
rect 296409 194147 296457 194175
rect 296485 194147 296519 194175
rect 296547 194147 296581 194175
rect 296609 194147 296643 194175
rect 296671 194147 296719 194175
rect 296409 194113 296719 194147
rect 296409 194085 296457 194113
rect 296485 194085 296519 194113
rect 296547 194085 296581 194113
rect 296609 194085 296643 194113
rect 296671 194085 296719 194113
rect 296409 194051 296719 194085
rect 296409 194023 296457 194051
rect 296485 194023 296519 194051
rect 296547 194023 296581 194051
rect 296609 194023 296643 194051
rect 296671 194023 296719 194051
rect 296409 193989 296719 194023
rect 296409 193961 296457 193989
rect 296485 193961 296519 193989
rect 296547 193961 296581 193989
rect 296609 193961 296643 193989
rect 296671 193961 296719 193989
rect 296409 185175 296719 193961
rect 296409 185147 296457 185175
rect 296485 185147 296519 185175
rect 296547 185147 296581 185175
rect 296609 185147 296643 185175
rect 296671 185147 296719 185175
rect 296409 185113 296719 185147
rect 296409 185085 296457 185113
rect 296485 185085 296519 185113
rect 296547 185085 296581 185113
rect 296609 185085 296643 185113
rect 296671 185085 296719 185113
rect 296409 185051 296719 185085
rect 296409 185023 296457 185051
rect 296485 185023 296519 185051
rect 296547 185023 296581 185051
rect 296609 185023 296643 185051
rect 296671 185023 296719 185051
rect 296409 184989 296719 185023
rect 296409 184961 296457 184989
rect 296485 184961 296519 184989
rect 296547 184961 296581 184989
rect 296609 184961 296643 184989
rect 296671 184961 296719 184989
rect 296409 176175 296719 184961
rect 296409 176147 296457 176175
rect 296485 176147 296519 176175
rect 296547 176147 296581 176175
rect 296609 176147 296643 176175
rect 296671 176147 296719 176175
rect 296409 176113 296719 176147
rect 296409 176085 296457 176113
rect 296485 176085 296519 176113
rect 296547 176085 296581 176113
rect 296609 176085 296643 176113
rect 296671 176085 296719 176113
rect 296409 176051 296719 176085
rect 296409 176023 296457 176051
rect 296485 176023 296519 176051
rect 296547 176023 296581 176051
rect 296609 176023 296643 176051
rect 296671 176023 296719 176051
rect 296409 175989 296719 176023
rect 296409 175961 296457 175989
rect 296485 175961 296519 175989
rect 296547 175961 296581 175989
rect 296609 175961 296643 175989
rect 296671 175961 296719 175989
rect 296409 167175 296719 175961
rect 296409 167147 296457 167175
rect 296485 167147 296519 167175
rect 296547 167147 296581 167175
rect 296609 167147 296643 167175
rect 296671 167147 296719 167175
rect 296409 167113 296719 167147
rect 296409 167085 296457 167113
rect 296485 167085 296519 167113
rect 296547 167085 296581 167113
rect 296609 167085 296643 167113
rect 296671 167085 296719 167113
rect 296409 167051 296719 167085
rect 296409 167023 296457 167051
rect 296485 167023 296519 167051
rect 296547 167023 296581 167051
rect 296609 167023 296643 167051
rect 296671 167023 296719 167051
rect 296409 166989 296719 167023
rect 296409 166961 296457 166989
rect 296485 166961 296519 166989
rect 296547 166961 296581 166989
rect 296609 166961 296643 166989
rect 296671 166961 296719 166989
rect 296409 158175 296719 166961
rect 296409 158147 296457 158175
rect 296485 158147 296519 158175
rect 296547 158147 296581 158175
rect 296609 158147 296643 158175
rect 296671 158147 296719 158175
rect 296409 158113 296719 158147
rect 296409 158085 296457 158113
rect 296485 158085 296519 158113
rect 296547 158085 296581 158113
rect 296609 158085 296643 158113
rect 296671 158085 296719 158113
rect 296409 158051 296719 158085
rect 296409 158023 296457 158051
rect 296485 158023 296519 158051
rect 296547 158023 296581 158051
rect 296609 158023 296643 158051
rect 296671 158023 296719 158051
rect 296409 157989 296719 158023
rect 296409 157961 296457 157989
rect 296485 157961 296519 157989
rect 296547 157961 296581 157989
rect 296609 157961 296643 157989
rect 296671 157961 296719 157989
rect 294549 146147 294597 146175
rect 294625 146147 294659 146175
rect 294687 146147 294721 146175
rect 294749 146147 294783 146175
rect 294811 146147 294859 146175
rect 294549 146113 294859 146147
rect 294549 146085 294597 146113
rect 294625 146085 294659 146113
rect 294687 146085 294721 146113
rect 294749 146085 294783 146113
rect 294811 146085 294859 146113
rect 294549 146051 294859 146085
rect 294549 146023 294597 146051
rect 294625 146023 294659 146051
rect 294687 146023 294721 146051
rect 294749 146023 294783 146051
rect 294811 146023 294859 146051
rect 294549 145989 294859 146023
rect 294549 145961 294597 145989
rect 294625 145961 294659 145989
rect 294687 145961 294721 145989
rect 294749 145961 294783 145989
rect 294811 145961 294859 145989
rect 294549 137175 294859 145961
rect 294549 137147 294597 137175
rect 294625 137147 294659 137175
rect 294687 137147 294721 137175
rect 294749 137147 294783 137175
rect 294811 137147 294859 137175
rect 294549 137113 294859 137147
rect 294549 137085 294597 137113
rect 294625 137085 294659 137113
rect 294687 137085 294721 137113
rect 294749 137085 294783 137113
rect 294811 137085 294859 137113
rect 294549 137051 294859 137085
rect 294549 137023 294597 137051
rect 294625 137023 294659 137051
rect 294687 137023 294721 137051
rect 294749 137023 294783 137051
rect 294811 137023 294859 137051
rect 294549 136989 294859 137023
rect 294549 136961 294597 136989
rect 294625 136961 294659 136989
rect 294687 136961 294721 136989
rect 294749 136961 294783 136989
rect 294811 136961 294859 136989
rect 294549 128175 294859 136961
rect 294549 128147 294597 128175
rect 294625 128147 294659 128175
rect 294687 128147 294721 128175
rect 294749 128147 294783 128175
rect 294811 128147 294859 128175
rect 294549 128113 294859 128147
rect 294549 128085 294597 128113
rect 294625 128085 294659 128113
rect 294687 128085 294721 128113
rect 294749 128085 294783 128113
rect 294811 128085 294859 128113
rect 294549 128051 294859 128085
rect 294549 128023 294597 128051
rect 294625 128023 294659 128051
rect 294687 128023 294721 128051
rect 294749 128023 294783 128051
rect 294811 128023 294859 128051
rect 294549 127989 294859 128023
rect 294549 127961 294597 127989
rect 294625 127961 294659 127989
rect 294687 127961 294721 127989
rect 294749 127961 294783 127989
rect 294811 127961 294859 127989
rect 294549 119175 294859 127961
rect 296409 149175 296719 157961
rect 296409 149147 296457 149175
rect 296485 149147 296519 149175
rect 296547 149147 296581 149175
rect 296609 149147 296643 149175
rect 296671 149147 296719 149175
rect 296409 149113 296719 149147
rect 296409 149085 296457 149113
rect 296485 149085 296519 149113
rect 296547 149085 296581 149113
rect 296609 149085 296643 149113
rect 296671 149085 296719 149113
rect 296409 149051 296719 149085
rect 296409 149023 296457 149051
rect 296485 149023 296519 149051
rect 296547 149023 296581 149051
rect 296609 149023 296643 149051
rect 296671 149023 296719 149051
rect 296409 148989 296719 149023
rect 296409 148961 296457 148989
rect 296485 148961 296519 148989
rect 296547 148961 296581 148989
rect 296609 148961 296643 148989
rect 296671 148961 296719 148989
rect 296409 140175 296719 148961
rect 296409 140147 296457 140175
rect 296485 140147 296519 140175
rect 296547 140147 296581 140175
rect 296609 140147 296643 140175
rect 296671 140147 296719 140175
rect 296409 140113 296719 140147
rect 296409 140085 296457 140113
rect 296485 140085 296519 140113
rect 296547 140085 296581 140113
rect 296609 140085 296643 140113
rect 296671 140085 296719 140113
rect 296409 140051 296719 140085
rect 296409 140023 296457 140051
rect 296485 140023 296519 140051
rect 296547 140023 296581 140051
rect 296609 140023 296643 140051
rect 296671 140023 296719 140051
rect 296409 139989 296719 140023
rect 296409 139961 296457 139989
rect 296485 139961 296519 139989
rect 296547 139961 296581 139989
rect 296609 139961 296643 139989
rect 296671 139961 296719 139989
rect 296409 131175 296719 139961
rect 296409 131147 296457 131175
rect 296485 131147 296519 131175
rect 296547 131147 296581 131175
rect 296609 131147 296643 131175
rect 296671 131147 296719 131175
rect 296409 131113 296719 131147
rect 296409 131085 296457 131113
rect 296485 131085 296519 131113
rect 296547 131085 296581 131113
rect 296609 131085 296643 131113
rect 296671 131085 296719 131113
rect 296409 131051 296719 131085
rect 296409 131023 296457 131051
rect 296485 131023 296519 131051
rect 296547 131023 296581 131051
rect 296609 131023 296643 131051
rect 296671 131023 296719 131051
rect 296409 130989 296719 131023
rect 296409 130961 296457 130989
rect 296485 130961 296519 130989
rect 296547 130961 296581 130989
rect 296609 130961 296643 130989
rect 296671 130961 296719 130989
rect 294549 119147 294597 119175
rect 294625 119147 294659 119175
rect 294687 119147 294721 119175
rect 294749 119147 294783 119175
rect 294811 119147 294859 119175
rect 294549 119113 294859 119147
rect 294549 119085 294597 119113
rect 294625 119085 294659 119113
rect 294687 119085 294721 119113
rect 294749 119085 294783 119113
rect 294811 119085 294859 119113
rect 294549 119051 294859 119085
rect 294549 119023 294597 119051
rect 294625 119023 294659 119051
rect 294687 119023 294721 119051
rect 294749 119023 294783 119051
rect 294811 119023 294859 119051
rect 294549 118989 294859 119023
rect 294549 118961 294597 118989
rect 294625 118961 294659 118989
rect 294687 118961 294721 118989
rect 294749 118961 294783 118989
rect 294811 118961 294859 118989
rect 294549 110175 294859 118961
rect 294549 110147 294597 110175
rect 294625 110147 294659 110175
rect 294687 110147 294721 110175
rect 294749 110147 294783 110175
rect 294811 110147 294859 110175
rect 294549 110113 294859 110147
rect 294549 110085 294597 110113
rect 294625 110085 294659 110113
rect 294687 110085 294721 110113
rect 294749 110085 294783 110113
rect 294811 110085 294859 110113
rect 294549 110051 294859 110085
rect 294549 110023 294597 110051
rect 294625 110023 294659 110051
rect 294687 110023 294721 110051
rect 294749 110023 294783 110051
rect 294811 110023 294859 110051
rect 294549 109989 294859 110023
rect 294549 109961 294597 109989
rect 294625 109961 294659 109989
rect 294687 109961 294721 109989
rect 294749 109961 294783 109989
rect 294811 109961 294859 109989
rect 294549 101175 294859 109961
rect 294549 101147 294597 101175
rect 294625 101147 294659 101175
rect 294687 101147 294721 101175
rect 294749 101147 294783 101175
rect 294811 101147 294859 101175
rect 294549 101113 294859 101147
rect 294549 101085 294597 101113
rect 294625 101085 294659 101113
rect 294687 101085 294721 101113
rect 294749 101085 294783 101113
rect 294811 101085 294859 101113
rect 294549 101051 294859 101085
rect 294549 101023 294597 101051
rect 294625 101023 294659 101051
rect 294687 101023 294721 101051
rect 294749 101023 294783 101051
rect 294811 101023 294859 101051
rect 294549 100989 294859 101023
rect 294549 100961 294597 100989
rect 294625 100961 294659 100989
rect 294687 100961 294721 100989
rect 294749 100961 294783 100989
rect 294811 100961 294859 100989
rect 294549 92175 294859 100961
rect 294549 92147 294597 92175
rect 294625 92147 294659 92175
rect 294687 92147 294721 92175
rect 294749 92147 294783 92175
rect 294811 92147 294859 92175
rect 294549 92113 294859 92147
rect 294549 92085 294597 92113
rect 294625 92085 294659 92113
rect 294687 92085 294721 92113
rect 294749 92085 294783 92113
rect 294811 92085 294859 92113
rect 294549 92051 294859 92085
rect 294549 92023 294597 92051
rect 294625 92023 294659 92051
rect 294687 92023 294721 92051
rect 294749 92023 294783 92051
rect 294811 92023 294859 92051
rect 294549 91989 294859 92023
rect 294549 91961 294597 91989
rect 294625 91961 294659 91989
rect 294687 91961 294721 91989
rect 294749 91961 294783 91989
rect 294811 91961 294859 91989
rect 294549 83175 294859 91961
rect 294549 83147 294597 83175
rect 294625 83147 294659 83175
rect 294687 83147 294721 83175
rect 294749 83147 294783 83175
rect 294811 83147 294859 83175
rect 294549 83113 294859 83147
rect 294549 83085 294597 83113
rect 294625 83085 294659 83113
rect 294687 83085 294721 83113
rect 294749 83085 294783 83113
rect 294811 83085 294859 83113
rect 294549 83051 294859 83085
rect 294549 83023 294597 83051
rect 294625 83023 294659 83051
rect 294687 83023 294721 83051
rect 294749 83023 294783 83051
rect 294811 83023 294859 83051
rect 294549 82989 294859 83023
rect 294549 82961 294597 82989
rect 294625 82961 294659 82989
rect 294687 82961 294721 82989
rect 294749 82961 294783 82989
rect 294811 82961 294859 82989
rect 294549 74175 294859 82961
rect 295246 125706 295274 125711
rect 295246 76370 295274 125678
rect 295358 125650 295386 125655
rect 295358 96194 295386 125622
rect 295470 125594 295498 125599
rect 295470 116018 295498 125566
rect 295470 115985 295498 115990
rect 296409 122175 296719 130961
rect 296409 122147 296457 122175
rect 296485 122147 296519 122175
rect 296547 122147 296581 122175
rect 296609 122147 296643 122175
rect 296671 122147 296719 122175
rect 296409 122113 296719 122147
rect 296409 122085 296457 122113
rect 296485 122085 296519 122113
rect 296547 122085 296581 122113
rect 296609 122085 296643 122113
rect 296671 122085 296719 122113
rect 296409 122051 296719 122085
rect 296409 122023 296457 122051
rect 296485 122023 296519 122051
rect 296547 122023 296581 122051
rect 296609 122023 296643 122051
rect 296671 122023 296719 122051
rect 296409 121989 296719 122023
rect 296409 121961 296457 121989
rect 296485 121961 296519 121989
rect 296547 121961 296581 121989
rect 296609 121961 296643 121989
rect 296671 121961 296719 121989
rect 295358 96161 295386 96166
rect 296409 113175 296719 121961
rect 296409 113147 296457 113175
rect 296485 113147 296519 113175
rect 296547 113147 296581 113175
rect 296609 113147 296643 113175
rect 296671 113147 296719 113175
rect 296409 113113 296719 113147
rect 296409 113085 296457 113113
rect 296485 113085 296519 113113
rect 296547 113085 296581 113113
rect 296609 113085 296643 113113
rect 296671 113085 296719 113113
rect 296409 113051 296719 113085
rect 296409 113023 296457 113051
rect 296485 113023 296519 113051
rect 296547 113023 296581 113051
rect 296609 113023 296643 113051
rect 296671 113023 296719 113051
rect 296409 112989 296719 113023
rect 296409 112961 296457 112989
rect 296485 112961 296519 112989
rect 296547 112961 296581 112989
rect 296609 112961 296643 112989
rect 296671 112961 296719 112989
rect 296409 104175 296719 112961
rect 296409 104147 296457 104175
rect 296485 104147 296519 104175
rect 296547 104147 296581 104175
rect 296609 104147 296643 104175
rect 296671 104147 296719 104175
rect 296409 104113 296719 104147
rect 296409 104085 296457 104113
rect 296485 104085 296519 104113
rect 296547 104085 296581 104113
rect 296609 104085 296643 104113
rect 296671 104085 296719 104113
rect 296409 104051 296719 104085
rect 296409 104023 296457 104051
rect 296485 104023 296519 104051
rect 296547 104023 296581 104051
rect 296609 104023 296643 104051
rect 296671 104023 296719 104051
rect 296409 103989 296719 104023
rect 296409 103961 296457 103989
rect 296485 103961 296519 103989
rect 296547 103961 296581 103989
rect 296609 103961 296643 103989
rect 296671 103961 296719 103989
rect 295246 76337 295274 76342
rect 296409 95175 296719 103961
rect 296409 95147 296457 95175
rect 296485 95147 296519 95175
rect 296547 95147 296581 95175
rect 296609 95147 296643 95175
rect 296671 95147 296719 95175
rect 296409 95113 296719 95147
rect 296409 95085 296457 95113
rect 296485 95085 296519 95113
rect 296547 95085 296581 95113
rect 296609 95085 296643 95113
rect 296671 95085 296719 95113
rect 296409 95051 296719 95085
rect 296409 95023 296457 95051
rect 296485 95023 296519 95051
rect 296547 95023 296581 95051
rect 296609 95023 296643 95051
rect 296671 95023 296719 95051
rect 296409 94989 296719 95023
rect 296409 94961 296457 94989
rect 296485 94961 296519 94989
rect 296547 94961 296581 94989
rect 296609 94961 296643 94989
rect 296671 94961 296719 94989
rect 296409 86175 296719 94961
rect 296409 86147 296457 86175
rect 296485 86147 296519 86175
rect 296547 86147 296581 86175
rect 296609 86147 296643 86175
rect 296671 86147 296719 86175
rect 296409 86113 296719 86147
rect 296409 86085 296457 86113
rect 296485 86085 296519 86113
rect 296547 86085 296581 86113
rect 296609 86085 296643 86113
rect 296671 86085 296719 86113
rect 296409 86051 296719 86085
rect 296409 86023 296457 86051
rect 296485 86023 296519 86051
rect 296547 86023 296581 86051
rect 296609 86023 296643 86051
rect 296671 86023 296719 86051
rect 296409 85989 296719 86023
rect 296409 85961 296457 85989
rect 296485 85961 296519 85989
rect 296547 85961 296581 85989
rect 296609 85961 296643 85989
rect 296671 85961 296719 85989
rect 296409 77175 296719 85961
rect 296409 77147 296457 77175
rect 296485 77147 296519 77175
rect 296547 77147 296581 77175
rect 296609 77147 296643 77175
rect 296671 77147 296719 77175
rect 296409 77113 296719 77147
rect 296409 77085 296457 77113
rect 296485 77085 296519 77113
rect 296547 77085 296581 77113
rect 296609 77085 296643 77113
rect 296671 77085 296719 77113
rect 296409 77051 296719 77085
rect 296409 77023 296457 77051
rect 296485 77023 296519 77051
rect 296547 77023 296581 77051
rect 296609 77023 296643 77051
rect 296671 77023 296719 77051
rect 296409 76989 296719 77023
rect 296409 76961 296457 76989
rect 296485 76961 296519 76989
rect 296547 76961 296581 76989
rect 296609 76961 296643 76989
rect 296671 76961 296719 76989
rect 294549 74147 294597 74175
rect 294625 74147 294659 74175
rect 294687 74147 294721 74175
rect 294749 74147 294783 74175
rect 294811 74147 294859 74175
rect 294549 74113 294859 74147
rect 294549 74085 294597 74113
rect 294625 74085 294659 74113
rect 294687 74085 294721 74113
rect 294749 74085 294783 74113
rect 294811 74085 294859 74113
rect 294549 74051 294859 74085
rect 294549 74023 294597 74051
rect 294625 74023 294659 74051
rect 294687 74023 294721 74051
rect 294749 74023 294783 74051
rect 294811 74023 294859 74051
rect 294549 73989 294859 74023
rect 294549 73961 294597 73989
rect 294625 73961 294659 73989
rect 294687 73961 294721 73989
rect 294749 73961 294783 73989
rect 294811 73961 294859 73989
rect 294549 65175 294859 73961
rect 294549 65147 294597 65175
rect 294625 65147 294659 65175
rect 294687 65147 294721 65175
rect 294749 65147 294783 65175
rect 294811 65147 294859 65175
rect 294549 65113 294859 65147
rect 294549 65085 294597 65113
rect 294625 65085 294659 65113
rect 294687 65085 294721 65113
rect 294749 65085 294783 65113
rect 294811 65085 294859 65113
rect 294549 65051 294859 65085
rect 294549 65023 294597 65051
rect 294625 65023 294659 65051
rect 294687 65023 294721 65051
rect 294749 65023 294783 65051
rect 294811 65023 294859 65051
rect 294549 64989 294859 65023
rect 294549 64961 294597 64989
rect 294625 64961 294659 64989
rect 294687 64961 294721 64989
rect 294749 64961 294783 64989
rect 294811 64961 294859 64989
rect 294549 56175 294859 64961
rect 294549 56147 294597 56175
rect 294625 56147 294659 56175
rect 294687 56147 294721 56175
rect 294749 56147 294783 56175
rect 294811 56147 294859 56175
rect 294549 56113 294859 56147
rect 294549 56085 294597 56113
rect 294625 56085 294659 56113
rect 294687 56085 294721 56113
rect 294749 56085 294783 56113
rect 294811 56085 294859 56113
rect 294549 56051 294859 56085
rect 294549 56023 294597 56051
rect 294625 56023 294659 56051
rect 294687 56023 294721 56051
rect 294749 56023 294783 56051
rect 294811 56023 294859 56051
rect 294549 55989 294859 56023
rect 294549 55961 294597 55989
rect 294625 55961 294659 55989
rect 294687 55961 294721 55989
rect 294749 55961 294783 55989
rect 294811 55961 294859 55989
rect 294549 47175 294859 55961
rect 294549 47147 294597 47175
rect 294625 47147 294659 47175
rect 294687 47147 294721 47175
rect 294749 47147 294783 47175
rect 294811 47147 294859 47175
rect 294549 47113 294859 47147
rect 294549 47085 294597 47113
rect 294625 47085 294659 47113
rect 294687 47085 294721 47113
rect 294749 47085 294783 47113
rect 294811 47085 294859 47113
rect 294549 47051 294859 47085
rect 294549 47023 294597 47051
rect 294625 47023 294659 47051
rect 294687 47023 294721 47051
rect 294749 47023 294783 47051
rect 294811 47023 294859 47051
rect 294549 46989 294859 47023
rect 294549 46961 294597 46989
rect 294625 46961 294659 46989
rect 294687 46961 294721 46989
rect 294749 46961 294783 46989
rect 294811 46961 294859 46989
rect 294549 38175 294859 46961
rect 294549 38147 294597 38175
rect 294625 38147 294659 38175
rect 294687 38147 294721 38175
rect 294749 38147 294783 38175
rect 294811 38147 294859 38175
rect 294549 38113 294859 38147
rect 294549 38085 294597 38113
rect 294625 38085 294659 38113
rect 294687 38085 294721 38113
rect 294749 38085 294783 38113
rect 294811 38085 294859 38113
rect 294549 38051 294859 38085
rect 294549 38023 294597 38051
rect 294625 38023 294659 38051
rect 294687 38023 294721 38051
rect 294749 38023 294783 38051
rect 294811 38023 294859 38051
rect 294549 37989 294859 38023
rect 294549 37961 294597 37989
rect 294625 37961 294659 37989
rect 294687 37961 294721 37989
rect 294749 37961 294783 37989
rect 294811 37961 294859 37989
rect 294549 29175 294859 37961
rect 294549 29147 294597 29175
rect 294625 29147 294659 29175
rect 294687 29147 294721 29175
rect 294749 29147 294783 29175
rect 294811 29147 294859 29175
rect 294549 29113 294859 29147
rect 294549 29085 294597 29113
rect 294625 29085 294659 29113
rect 294687 29085 294721 29113
rect 294749 29085 294783 29113
rect 294811 29085 294859 29113
rect 294549 29051 294859 29085
rect 294549 29023 294597 29051
rect 294625 29023 294659 29051
rect 294687 29023 294721 29051
rect 294749 29023 294783 29051
rect 294811 29023 294859 29051
rect 294549 28989 294859 29023
rect 294549 28961 294597 28989
rect 294625 28961 294659 28989
rect 294687 28961 294721 28989
rect 294749 28961 294783 28989
rect 294811 28961 294859 28989
rect 294549 20175 294859 28961
rect 294549 20147 294597 20175
rect 294625 20147 294659 20175
rect 294687 20147 294721 20175
rect 294749 20147 294783 20175
rect 294811 20147 294859 20175
rect 294549 20113 294859 20147
rect 294549 20085 294597 20113
rect 294625 20085 294659 20113
rect 294687 20085 294721 20113
rect 294749 20085 294783 20113
rect 294811 20085 294859 20113
rect 294549 20051 294859 20085
rect 294549 20023 294597 20051
rect 294625 20023 294659 20051
rect 294687 20023 294721 20051
rect 294749 20023 294783 20051
rect 294811 20023 294859 20051
rect 294549 19989 294859 20023
rect 294549 19961 294597 19989
rect 294625 19961 294659 19989
rect 294687 19961 294721 19989
rect 294749 19961 294783 19989
rect 294811 19961 294859 19989
rect 294549 11175 294859 19961
rect 294549 11147 294597 11175
rect 294625 11147 294659 11175
rect 294687 11147 294721 11175
rect 294749 11147 294783 11175
rect 294811 11147 294859 11175
rect 294549 11113 294859 11147
rect 294549 11085 294597 11113
rect 294625 11085 294659 11113
rect 294687 11085 294721 11113
rect 294749 11085 294783 11113
rect 294811 11085 294859 11113
rect 294549 11051 294859 11085
rect 294549 11023 294597 11051
rect 294625 11023 294659 11051
rect 294687 11023 294721 11051
rect 294749 11023 294783 11051
rect 294811 11023 294859 11051
rect 294549 10989 294859 11023
rect 294549 10961 294597 10989
rect 294625 10961 294659 10989
rect 294687 10961 294721 10989
rect 294749 10961 294783 10989
rect 294811 10961 294859 10989
rect 294549 2175 294859 10961
rect 294549 2147 294597 2175
rect 294625 2147 294659 2175
rect 294687 2147 294721 2175
rect 294749 2147 294783 2175
rect 294811 2147 294859 2175
rect 294549 2113 294859 2147
rect 294549 2085 294597 2113
rect 294625 2085 294659 2113
rect 294687 2085 294721 2113
rect 294749 2085 294783 2113
rect 294811 2085 294859 2113
rect 294549 2051 294859 2085
rect 294549 2023 294597 2051
rect 294625 2023 294659 2051
rect 294687 2023 294721 2051
rect 294749 2023 294783 2051
rect 294811 2023 294859 2051
rect 294549 1989 294859 2023
rect 294549 1961 294597 1989
rect 294625 1961 294659 1989
rect 294687 1961 294721 1989
rect 294749 1961 294783 1989
rect 294811 1961 294859 1989
rect 294549 -80 294859 1961
rect 294549 -108 294597 -80
rect 294625 -108 294659 -80
rect 294687 -108 294721 -80
rect 294749 -108 294783 -80
rect 294811 -108 294859 -80
rect 294549 -142 294859 -108
rect 294549 -170 294597 -142
rect 294625 -170 294659 -142
rect 294687 -170 294721 -142
rect 294749 -170 294783 -142
rect 294811 -170 294859 -142
rect 294549 -204 294859 -170
rect 294549 -232 294597 -204
rect 294625 -232 294659 -204
rect 294687 -232 294721 -204
rect 294749 -232 294783 -204
rect 294811 -232 294859 -204
rect 294549 -266 294859 -232
rect 294549 -294 294597 -266
rect 294625 -294 294659 -266
rect 294687 -294 294721 -266
rect 294749 -294 294783 -266
rect 294811 -294 294859 -266
rect 294549 -822 294859 -294
rect 296409 68175 296719 76961
rect 296409 68147 296457 68175
rect 296485 68147 296519 68175
rect 296547 68147 296581 68175
rect 296609 68147 296643 68175
rect 296671 68147 296719 68175
rect 296409 68113 296719 68147
rect 296409 68085 296457 68113
rect 296485 68085 296519 68113
rect 296547 68085 296581 68113
rect 296609 68085 296643 68113
rect 296671 68085 296719 68113
rect 296409 68051 296719 68085
rect 296409 68023 296457 68051
rect 296485 68023 296519 68051
rect 296547 68023 296581 68051
rect 296609 68023 296643 68051
rect 296671 68023 296719 68051
rect 296409 67989 296719 68023
rect 296409 67961 296457 67989
rect 296485 67961 296519 67989
rect 296547 67961 296581 67989
rect 296609 67961 296643 67989
rect 296671 67961 296719 67989
rect 296409 59175 296719 67961
rect 296409 59147 296457 59175
rect 296485 59147 296519 59175
rect 296547 59147 296581 59175
rect 296609 59147 296643 59175
rect 296671 59147 296719 59175
rect 296409 59113 296719 59147
rect 296409 59085 296457 59113
rect 296485 59085 296519 59113
rect 296547 59085 296581 59113
rect 296609 59085 296643 59113
rect 296671 59085 296719 59113
rect 296409 59051 296719 59085
rect 296409 59023 296457 59051
rect 296485 59023 296519 59051
rect 296547 59023 296581 59051
rect 296609 59023 296643 59051
rect 296671 59023 296719 59051
rect 296409 58989 296719 59023
rect 296409 58961 296457 58989
rect 296485 58961 296519 58989
rect 296547 58961 296581 58989
rect 296609 58961 296643 58989
rect 296671 58961 296719 58989
rect 296409 50175 296719 58961
rect 296409 50147 296457 50175
rect 296485 50147 296519 50175
rect 296547 50147 296581 50175
rect 296609 50147 296643 50175
rect 296671 50147 296719 50175
rect 296409 50113 296719 50147
rect 296409 50085 296457 50113
rect 296485 50085 296519 50113
rect 296547 50085 296581 50113
rect 296609 50085 296643 50113
rect 296671 50085 296719 50113
rect 296409 50051 296719 50085
rect 296409 50023 296457 50051
rect 296485 50023 296519 50051
rect 296547 50023 296581 50051
rect 296609 50023 296643 50051
rect 296671 50023 296719 50051
rect 296409 49989 296719 50023
rect 296409 49961 296457 49989
rect 296485 49961 296519 49989
rect 296547 49961 296581 49989
rect 296609 49961 296643 49989
rect 296671 49961 296719 49989
rect 296409 41175 296719 49961
rect 296409 41147 296457 41175
rect 296485 41147 296519 41175
rect 296547 41147 296581 41175
rect 296609 41147 296643 41175
rect 296671 41147 296719 41175
rect 296409 41113 296719 41147
rect 296409 41085 296457 41113
rect 296485 41085 296519 41113
rect 296547 41085 296581 41113
rect 296609 41085 296643 41113
rect 296671 41085 296719 41113
rect 296409 41051 296719 41085
rect 296409 41023 296457 41051
rect 296485 41023 296519 41051
rect 296547 41023 296581 41051
rect 296609 41023 296643 41051
rect 296671 41023 296719 41051
rect 296409 40989 296719 41023
rect 296409 40961 296457 40989
rect 296485 40961 296519 40989
rect 296547 40961 296581 40989
rect 296609 40961 296643 40989
rect 296671 40961 296719 40989
rect 296409 32175 296719 40961
rect 296409 32147 296457 32175
rect 296485 32147 296519 32175
rect 296547 32147 296581 32175
rect 296609 32147 296643 32175
rect 296671 32147 296719 32175
rect 296409 32113 296719 32147
rect 296409 32085 296457 32113
rect 296485 32085 296519 32113
rect 296547 32085 296581 32113
rect 296609 32085 296643 32113
rect 296671 32085 296719 32113
rect 296409 32051 296719 32085
rect 296409 32023 296457 32051
rect 296485 32023 296519 32051
rect 296547 32023 296581 32051
rect 296609 32023 296643 32051
rect 296671 32023 296719 32051
rect 296409 31989 296719 32023
rect 296409 31961 296457 31989
rect 296485 31961 296519 31989
rect 296547 31961 296581 31989
rect 296609 31961 296643 31989
rect 296671 31961 296719 31989
rect 296409 23175 296719 31961
rect 296409 23147 296457 23175
rect 296485 23147 296519 23175
rect 296547 23147 296581 23175
rect 296609 23147 296643 23175
rect 296671 23147 296719 23175
rect 296409 23113 296719 23147
rect 296409 23085 296457 23113
rect 296485 23085 296519 23113
rect 296547 23085 296581 23113
rect 296609 23085 296643 23113
rect 296671 23085 296719 23113
rect 296409 23051 296719 23085
rect 296409 23023 296457 23051
rect 296485 23023 296519 23051
rect 296547 23023 296581 23051
rect 296609 23023 296643 23051
rect 296671 23023 296719 23051
rect 296409 22989 296719 23023
rect 296409 22961 296457 22989
rect 296485 22961 296519 22989
rect 296547 22961 296581 22989
rect 296609 22961 296643 22989
rect 296671 22961 296719 22989
rect 296409 14175 296719 22961
rect 296409 14147 296457 14175
rect 296485 14147 296519 14175
rect 296547 14147 296581 14175
rect 296609 14147 296643 14175
rect 296671 14147 296719 14175
rect 296409 14113 296719 14147
rect 296409 14085 296457 14113
rect 296485 14085 296519 14113
rect 296547 14085 296581 14113
rect 296609 14085 296643 14113
rect 296671 14085 296719 14113
rect 296409 14051 296719 14085
rect 296409 14023 296457 14051
rect 296485 14023 296519 14051
rect 296547 14023 296581 14051
rect 296609 14023 296643 14051
rect 296671 14023 296719 14051
rect 296409 13989 296719 14023
rect 296409 13961 296457 13989
rect 296485 13961 296519 13989
rect 296547 13961 296581 13989
rect 296609 13961 296643 13989
rect 296671 13961 296719 13989
rect 296409 5175 296719 13961
rect 296409 5147 296457 5175
rect 296485 5147 296519 5175
rect 296547 5147 296581 5175
rect 296609 5147 296643 5175
rect 296671 5147 296719 5175
rect 296409 5113 296719 5147
rect 296409 5085 296457 5113
rect 296485 5085 296519 5113
rect 296547 5085 296581 5113
rect 296609 5085 296643 5113
rect 296671 5085 296719 5113
rect 296409 5051 296719 5085
rect 296409 5023 296457 5051
rect 296485 5023 296519 5051
rect 296547 5023 296581 5051
rect 296609 5023 296643 5051
rect 296671 5023 296719 5051
rect 296409 4989 296719 5023
rect 296409 4961 296457 4989
rect 296485 4961 296519 4989
rect 296547 4961 296581 4989
rect 296609 4961 296643 4989
rect 296671 4961 296719 4989
rect 296409 -560 296719 4961
rect 298200 298606 298510 298654
rect 298200 298578 298248 298606
rect 298276 298578 298310 298606
rect 298338 298578 298372 298606
rect 298400 298578 298434 298606
rect 298462 298578 298510 298606
rect 298200 298544 298510 298578
rect 298200 298516 298248 298544
rect 298276 298516 298310 298544
rect 298338 298516 298372 298544
rect 298400 298516 298434 298544
rect 298462 298516 298510 298544
rect 298200 298482 298510 298516
rect 298200 298454 298248 298482
rect 298276 298454 298310 298482
rect 298338 298454 298372 298482
rect 298400 298454 298434 298482
rect 298462 298454 298510 298482
rect 298200 298420 298510 298454
rect 298200 298392 298248 298420
rect 298276 298392 298310 298420
rect 298338 298392 298372 298420
rect 298400 298392 298434 298420
rect 298462 298392 298510 298420
rect 298200 290175 298510 298392
rect 298200 290147 298248 290175
rect 298276 290147 298310 290175
rect 298338 290147 298372 290175
rect 298400 290147 298434 290175
rect 298462 290147 298510 290175
rect 298200 290113 298510 290147
rect 298200 290085 298248 290113
rect 298276 290085 298310 290113
rect 298338 290085 298372 290113
rect 298400 290085 298434 290113
rect 298462 290085 298510 290113
rect 298200 290051 298510 290085
rect 298200 290023 298248 290051
rect 298276 290023 298310 290051
rect 298338 290023 298372 290051
rect 298400 290023 298434 290051
rect 298462 290023 298510 290051
rect 298200 289989 298510 290023
rect 298200 289961 298248 289989
rect 298276 289961 298310 289989
rect 298338 289961 298372 289989
rect 298400 289961 298434 289989
rect 298462 289961 298510 289989
rect 298200 281175 298510 289961
rect 298200 281147 298248 281175
rect 298276 281147 298310 281175
rect 298338 281147 298372 281175
rect 298400 281147 298434 281175
rect 298462 281147 298510 281175
rect 298200 281113 298510 281147
rect 298200 281085 298248 281113
rect 298276 281085 298310 281113
rect 298338 281085 298372 281113
rect 298400 281085 298434 281113
rect 298462 281085 298510 281113
rect 298200 281051 298510 281085
rect 298200 281023 298248 281051
rect 298276 281023 298310 281051
rect 298338 281023 298372 281051
rect 298400 281023 298434 281051
rect 298462 281023 298510 281051
rect 298200 280989 298510 281023
rect 298200 280961 298248 280989
rect 298276 280961 298310 280989
rect 298338 280961 298372 280989
rect 298400 280961 298434 280989
rect 298462 280961 298510 280989
rect 298200 272175 298510 280961
rect 298200 272147 298248 272175
rect 298276 272147 298310 272175
rect 298338 272147 298372 272175
rect 298400 272147 298434 272175
rect 298462 272147 298510 272175
rect 298200 272113 298510 272147
rect 298200 272085 298248 272113
rect 298276 272085 298310 272113
rect 298338 272085 298372 272113
rect 298400 272085 298434 272113
rect 298462 272085 298510 272113
rect 298200 272051 298510 272085
rect 298200 272023 298248 272051
rect 298276 272023 298310 272051
rect 298338 272023 298372 272051
rect 298400 272023 298434 272051
rect 298462 272023 298510 272051
rect 298200 271989 298510 272023
rect 298200 271961 298248 271989
rect 298276 271961 298310 271989
rect 298338 271961 298372 271989
rect 298400 271961 298434 271989
rect 298462 271961 298510 271989
rect 298200 263175 298510 271961
rect 298200 263147 298248 263175
rect 298276 263147 298310 263175
rect 298338 263147 298372 263175
rect 298400 263147 298434 263175
rect 298462 263147 298510 263175
rect 298200 263113 298510 263147
rect 298200 263085 298248 263113
rect 298276 263085 298310 263113
rect 298338 263085 298372 263113
rect 298400 263085 298434 263113
rect 298462 263085 298510 263113
rect 298200 263051 298510 263085
rect 298200 263023 298248 263051
rect 298276 263023 298310 263051
rect 298338 263023 298372 263051
rect 298400 263023 298434 263051
rect 298462 263023 298510 263051
rect 298200 262989 298510 263023
rect 298200 262961 298248 262989
rect 298276 262961 298310 262989
rect 298338 262961 298372 262989
rect 298400 262961 298434 262989
rect 298462 262961 298510 262989
rect 298200 254175 298510 262961
rect 298200 254147 298248 254175
rect 298276 254147 298310 254175
rect 298338 254147 298372 254175
rect 298400 254147 298434 254175
rect 298462 254147 298510 254175
rect 298200 254113 298510 254147
rect 298200 254085 298248 254113
rect 298276 254085 298310 254113
rect 298338 254085 298372 254113
rect 298400 254085 298434 254113
rect 298462 254085 298510 254113
rect 298200 254051 298510 254085
rect 298200 254023 298248 254051
rect 298276 254023 298310 254051
rect 298338 254023 298372 254051
rect 298400 254023 298434 254051
rect 298462 254023 298510 254051
rect 298200 253989 298510 254023
rect 298200 253961 298248 253989
rect 298276 253961 298310 253989
rect 298338 253961 298372 253989
rect 298400 253961 298434 253989
rect 298462 253961 298510 253989
rect 298200 245175 298510 253961
rect 298200 245147 298248 245175
rect 298276 245147 298310 245175
rect 298338 245147 298372 245175
rect 298400 245147 298434 245175
rect 298462 245147 298510 245175
rect 298200 245113 298510 245147
rect 298200 245085 298248 245113
rect 298276 245085 298310 245113
rect 298338 245085 298372 245113
rect 298400 245085 298434 245113
rect 298462 245085 298510 245113
rect 298200 245051 298510 245085
rect 298200 245023 298248 245051
rect 298276 245023 298310 245051
rect 298338 245023 298372 245051
rect 298400 245023 298434 245051
rect 298462 245023 298510 245051
rect 298200 244989 298510 245023
rect 298200 244961 298248 244989
rect 298276 244961 298310 244989
rect 298338 244961 298372 244989
rect 298400 244961 298434 244989
rect 298462 244961 298510 244989
rect 298200 236175 298510 244961
rect 298200 236147 298248 236175
rect 298276 236147 298310 236175
rect 298338 236147 298372 236175
rect 298400 236147 298434 236175
rect 298462 236147 298510 236175
rect 298200 236113 298510 236147
rect 298200 236085 298248 236113
rect 298276 236085 298310 236113
rect 298338 236085 298372 236113
rect 298400 236085 298434 236113
rect 298462 236085 298510 236113
rect 298200 236051 298510 236085
rect 298200 236023 298248 236051
rect 298276 236023 298310 236051
rect 298338 236023 298372 236051
rect 298400 236023 298434 236051
rect 298462 236023 298510 236051
rect 298200 235989 298510 236023
rect 298200 235961 298248 235989
rect 298276 235961 298310 235989
rect 298338 235961 298372 235989
rect 298400 235961 298434 235989
rect 298462 235961 298510 235989
rect 298200 227175 298510 235961
rect 298200 227147 298248 227175
rect 298276 227147 298310 227175
rect 298338 227147 298372 227175
rect 298400 227147 298434 227175
rect 298462 227147 298510 227175
rect 298200 227113 298510 227147
rect 298200 227085 298248 227113
rect 298276 227085 298310 227113
rect 298338 227085 298372 227113
rect 298400 227085 298434 227113
rect 298462 227085 298510 227113
rect 298200 227051 298510 227085
rect 298200 227023 298248 227051
rect 298276 227023 298310 227051
rect 298338 227023 298372 227051
rect 298400 227023 298434 227051
rect 298462 227023 298510 227051
rect 298200 226989 298510 227023
rect 298200 226961 298248 226989
rect 298276 226961 298310 226989
rect 298338 226961 298372 226989
rect 298400 226961 298434 226989
rect 298462 226961 298510 226989
rect 298200 218175 298510 226961
rect 298200 218147 298248 218175
rect 298276 218147 298310 218175
rect 298338 218147 298372 218175
rect 298400 218147 298434 218175
rect 298462 218147 298510 218175
rect 298200 218113 298510 218147
rect 298200 218085 298248 218113
rect 298276 218085 298310 218113
rect 298338 218085 298372 218113
rect 298400 218085 298434 218113
rect 298462 218085 298510 218113
rect 298200 218051 298510 218085
rect 298200 218023 298248 218051
rect 298276 218023 298310 218051
rect 298338 218023 298372 218051
rect 298400 218023 298434 218051
rect 298462 218023 298510 218051
rect 298200 217989 298510 218023
rect 298200 217961 298248 217989
rect 298276 217961 298310 217989
rect 298338 217961 298372 217989
rect 298400 217961 298434 217989
rect 298462 217961 298510 217989
rect 298200 209175 298510 217961
rect 298200 209147 298248 209175
rect 298276 209147 298310 209175
rect 298338 209147 298372 209175
rect 298400 209147 298434 209175
rect 298462 209147 298510 209175
rect 298200 209113 298510 209147
rect 298200 209085 298248 209113
rect 298276 209085 298310 209113
rect 298338 209085 298372 209113
rect 298400 209085 298434 209113
rect 298462 209085 298510 209113
rect 298200 209051 298510 209085
rect 298200 209023 298248 209051
rect 298276 209023 298310 209051
rect 298338 209023 298372 209051
rect 298400 209023 298434 209051
rect 298462 209023 298510 209051
rect 298200 208989 298510 209023
rect 298200 208961 298248 208989
rect 298276 208961 298310 208989
rect 298338 208961 298372 208989
rect 298400 208961 298434 208989
rect 298462 208961 298510 208989
rect 298200 200175 298510 208961
rect 298200 200147 298248 200175
rect 298276 200147 298310 200175
rect 298338 200147 298372 200175
rect 298400 200147 298434 200175
rect 298462 200147 298510 200175
rect 298200 200113 298510 200147
rect 298200 200085 298248 200113
rect 298276 200085 298310 200113
rect 298338 200085 298372 200113
rect 298400 200085 298434 200113
rect 298462 200085 298510 200113
rect 298200 200051 298510 200085
rect 298200 200023 298248 200051
rect 298276 200023 298310 200051
rect 298338 200023 298372 200051
rect 298400 200023 298434 200051
rect 298462 200023 298510 200051
rect 298200 199989 298510 200023
rect 298200 199961 298248 199989
rect 298276 199961 298310 199989
rect 298338 199961 298372 199989
rect 298400 199961 298434 199989
rect 298462 199961 298510 199989
rect 298200 191175 298510 199961
rect 298200 191147 298248 191175
rect 298276 191147 298310 191175
rect 298338 191147 298372 191175
rect 298400 191147 298434 191175
rect 298462 191147 298510 191175
rect 298200 191113 298510 191147
rect 298200 191085 298248 191113
rect 298276 191085 298310 191113
rect 298338 191085 298372 191113
rect 298400 191085 298434 191113
rect 298462 191085 298510 191113
rect 298200 191051 298510 191085
rect 298200 191023 298248 191051
rect 298276 191023 298310 191051
rect 298338 191023 298372 191051
rect 298400 191023 298434 191051
rect 298462 191023 298510 191051
rect 298200 190989 298510 191023
rect 298200 190961 298248 190989
rect 298276 190961 298310 190989
rect 298338 190961 298372 190989
rect 298400 190961 298434 190989
rect 298462 190961 298510 190989
rect 298200 182175 298510 190961
rect 298200 182147 298248 182175
rect 298276 182147 298310 182175
rect 298338 182147 298372 182175
rect 298400 182147 298434 182175
rect 298462 182147 298510 182175
rect 298200 182113 298510 182147
rect 298200 182085 298248 182113
rect 298276 182085 298310 182113
rect 298338 182085 298372 182113
rect 298400 182085 298434 182113
rect 298462 182085 298510 182113
rect 298200 182051 298510 182085
rect 298200 182023 298248 182051
rect 298276 182023 298310 182051
rect 298338 182023 298372 182051
rect 298400 182023 298434 182051
rect 298462 182023 298510 182051
rect 298200 181989 298510 182023
rect 298200 181961 298248 181989
rect 298276 181961 298310 181989
rect 298338 181961 298372 181989
rect 298400 181961 298434 181989
rect 298462 181961 298510 181989
rect 298200 173175 298510 181961
rect 298200 173147 298248 173175
rect 298276 173147 298310 173175
rect 298338 173147 298372 173175
rect 298400 173147 298434 173175
rect 298462 173147 298510 173175
rect 298200 173113 298510 173147
rect 298200 173085 298248 173113
rect 298276 173085 298310 173113
rect 298338 173085 298372 173113
rect 298400 173085 298434 173113
rect 298462 173085 298510 173113
rect 298200 173051 298510 173085
rect 298200 173023 298248 173051
rect 298276 173023 298310 173051
rect 298338 173023 298372 173051
rect 298400 173023 298434 173051
rect 298462 173023 298510 173051
rect 298200 172989 298510 173023
rect 298200 172961 298248 172989
rect 298276 172961 298310 172989
rect 298338 172961 298372 172989
rect 298400 172961 298434 172989
rect 298462 172961 298510 172989
rect 298200 164175 298510 172961
rect 298200 164147 298248 164175
rect 298276 164147 298310 164175
rect 298338 164147 298372 164175
rect 298400 164147 298434 164175
rect 298462 164147 298510 164175
rect 298200 164113 298510 164147
rect 298200 164085 298248 164113
rect 298276 164085 298310 164113
rect 298338 164085 298372 164113
rect 298400 164085 298434 164113
rect 298462 164085 298510 164113
rect 298200 164051 298510 164085
rect 298200 164023 298248 164051
rect 298276 164023 298310 164051
rect 298338 164023 298372 164051
rect 298400 164023 298434 164051
rect 298462 164023 298510 164051
rect 298200 163989 298510 164023
rect 298200 163961 298248 163989
rect 298276 163961 298310 163989
rect 298338 163961 298372 163989
rect 298400 163961 298434 163989
rect 298462 163961 298510 163989
rect 298200 155175 298510 163961
rect 298200 155147 298248 155175
rect 298276 155147 298310 155175
rect 298338 155147 298372 155175
rect 298400 155147 298434 155175
rect 298462 155147 298510 155175
rect 298200 155113 298510 155147
rect 298200 155085 298248 155113
rect 298276 155085 298310 155113
rect 298338 155085 298372 155113
rect 298400 155085 298434 155113
rect 298462 155085 298510 155113
rect 298200 155051 298510 155085
rect 298200 155023 298248 155051
rect 298276 155023 298310 155051
rect 298338 155023 298372 155051
rect 298400 155023 298434 155051
rect 298462 155023 298510 155051
rect 298200 154989 298510 155023
rect 298200 154961 298248 154989
rect 298276 154961 298310 154989
rect 298338 154961 298372 154989
rect 298400 154961 298434 154989
rect 298462 154961 298510 154989
rect 298200 146175 298510 154961
rect 298200 146147 298248 146175
rect 298276 146147 298310 146175
rect 298338 146147 298372 146175
rect 298400 146147 298434 146175
rect 298462 146147 298510 146175
rect 298200 146113 298510 146147
rect 298200 146085 298248 146113
rect 298276 146085 298310 146113
rect 298338 146085 298372 146113
rect 298400 146085 298434 146113
rect 298462 146085 298510 146113
rect 298200 146051 298510 146085
rect 298200 146023 298248 146051
rect 298276 146023 298310 146051
rect 298338 146023 298372 146051
rect 298400 146023 298434 146051
rect 298462 146023 298510 146051
rect 298200 145989 298510 146023
rect 298200 145961 298248 145989
rect 298276 145961 298310 145989
rect 298338 145961 298372 145989
rect 298400 145961 298434 145989
rect 298462 145961 298510 145989
rect 298200 137175 298510 145961
rect 298200 137147 298248 137175
rect 298276 137147 298310 137175
rect 298338 137147 298372 137175
rect 298400 137147 298434 137175
rect 298462 137147 298510 137175
rect 298200 137113 298510 137147
rect 298200 137085 298248 137113
rect 298276 137085 298310 137113
rect 298338 137085 298372 137113
rect 298400 137085 298434 137113
rect 298462 137085 298510 137113
rect 298200 137051 298510 137085
rect 298200 137023 298248 137051
rect 298276 137023 298310 137051
rect 298338 137023 298372 137051
rect 298400 137023 298434 137051
rect 298462 137023 298510 137051
rect 298200 136989 298510 137023
rect 298200 136961 298248 136989
rect 298276 136961 298310 136989
rect 298338 136961 298372 136989
rect 298400 136961 298434 136989
rect 298462 136961 298510 136989
rect 298200 128175 298510 136961
rect 298200 128147 298248 128175
rect 298276 128147 298310 128175
rect 298338 128147 298372 128175
rect 298400 128147 298434 128175
rect 298462 128147 298510 128175
rect 298200 128113 298510 128147
rect 298200 128085 298248 128113
rect 298276 128085 298310 128113
rect 298338 128085 298372 128113
rect 298400 128085 298434 128113
rect 298462 128085 298510 128113
rect 298200 128051 298510 128085
rect 298200 128023 298248 128051
rect 298276 128023 298310 128051
rect 298338 128023 298372 128051
rect 298400 128023 298434 128051
rect 298462 128023 298510 128051
rect 298200 127989 298510 128023
rect 298200 127961 298248 127989
rect 298276 127961 298310 127989
rect 298338 127961 298372 127989
rect 298400 127961 298434 127989
rect 298462 127961 298510 127989
rect 298200 119175 298510 127961
rect 298200 119147 298248 119175
rect 298276 119147 298310 119175
rect 298338 119147 298372 119175
rect 298400 119147 298434 119175
rect 298462 119147 298510 119175
rect 298200 119113 298510 119147
rect 298200 119085 298248 119113
rect 298276 119085 298310 119113
rect 298338 119085 298372 119113
rect 298400 119085 298434 119113
rect 298462 119085 298510 119113
rect 298200 119051 298510 119085
rect 298200 119023 298248 119051
rect 298276 119023 298310 119051
rect 298338 119023 298372 119051
rect 298400 119023 298434 119051
rect 298462 119023 298510 119051
rect 298200 118989 298510 119023
rect 298200 118961 298248 118989
rect 298276 118961 298310 118989
rect 298338 118961 298372 118989
rect 298400 118961 298434 118989
rect 298462 118961 298510 118989
rect 298200 110175 298510 118961
rect 298200 110147 298248 110175
rect 298276 110147 298310 110175
rect 298338 110147 298372 110175
rect 298400 110147 298434 110175
rect 298462 110147 298510 110175
rect 298200 110113 298510 110147
rect 298200 110085 298248 110113
rect 298276 110085 298310 110113
rect 298338 110085 298372 110113
rect 298400 110085 298434 110113
rect 298462 110085 298510 110113
rect 298200 110051 298510 110085
rect 298200 110023 298248 110051
rect 298276 110023 298310 110051
rect 298338 110023 298372 110051
rect 298400 110023 298434 110051
rect 298462 110023 298510 110051
rect 298200 109989 298510 110023
rect 298200 109961 298248 109989
rect 298276 109961 298310 109989
rect 298338 109961 298372 109989
rect 298400 109961 298434 109989
rect 298462 109961 298510 109989
rect 298200 101175 298510 109961
rect 298200 101147 298248 101175
rect 298276 101147 298310 101175
rect 298338 101147 298372 101175
rect 298400 101147 298434 101175
rect 298462 101147 298510 101175
rect 298200 101113 298510 101147
rect 298200 101085 298248 101113
rect 298276 101085 298310 101113
rect 298338 101085 298372 101113
rect 298400 101085 298434 101113
rect 298462 101085 298510 101113
rect 298200 101051 298510 101085
rect 298200 101023 298248 101051
rect 298276 101023 298310 101051
rect 298338 101023 298372 101051
rect 298400 101023 298434 101051
rect 298462 101023 298510 101051
rect 298200 100989 298510 101023
rect 298200 100961 298248 100989
rect 298276 100961 298310 100989
rect 298338 100961 298372 100989
rect 298400 100961 298434 100989
rect 298462 100961 298510 100989
rect 298200 92175 298510 100961
rect 298200 92147 298248 92175
rect 298276 92147 298310 92175
rect 298338 92147 298372 92175
rect 298400 92147 298434 92175
rect 298462 92147 298510 92175
rect 298200 92113 298510 92147
rect 298200 92085 298248 92113
rect 298276 92085 298310 92113
rect 298338 92085 298372 92113
rect 298400 92085 298434 92113
rect 298462 92085 298510 92113
rect 298200 92051 298510 92085
rect 298200 92023 298248 92051
rect 298276 92023 298310 92051
rect 298338 92023 298372 92051
rect 298400 92023 298434 92051
rect 298462 92023 298510 92051
rect 298200 91989 298510 92023
rect 298200 91961 298248 91989
rect 298276 91961 298310 91989
rect 298338 91961 298372 91989
rect 298400 91961 298434 91989
rect 298462 91961 298510 91989
rect 298200 83175 298510 91961
rect 298200 83147 298248 83175
rect 298276 83147 298310 83175
rect 298338 83147 298372 83175
rect 298400 83147 298434 83175
rect 298462 83147 298510 83175
rect 298200 83113 298510 83147
rect 298200 83085 298248 83113
rect 298276 83085 298310 83113
rect 298338 83085 298372 83113
rect 298400 83085 298434 83113
rect 298462 83085 298510 83113
rect 298200 83051 298510 83085
rect 298200 83023 298248 83051
rect 298276 83023 298310 83051
rect 298338 83023 298372 83051
rect 298400 83023 298434 83051
rect 298462 83023 298510 83051
rect 298200 82989 298510 83023
rect 298200 82961 298248 82989
rect 298276 82961 298310 82989
rect 298338 82961 298372 82989
rect 298400 82961 298434 82989
rect 298462 82961 298510 82989
rect 298200 74175 298510 82961
rect 298200 74147 298248 74175
rect 298276 74147 298310 74175
rect 298338 74147 298372 74175
rect 298400 74147 298434 74175
rect 298462 74147 298510 74175
rect 298200 74113 298510 74147
rect 298200 74085 298248 74113
rect 298276 74085 298310 74113
rect 298338 74085 298372 74113
rect 298400 74085 298434 74113
rect 298462 74085 298510 74113
rect 298200 74051 298510 74085
rect 298200 74023 298248 74051
rect 298276 74023 298310 74051
rect 298338 74023 298372 74051
rect 298400 74023 298434 74051
rect 298462 74023 298510 74051
rect 298200 73989 298510 74023
rect 298200 73961 298248 73989
rect 298276 73961 298310 73989
rect 298338 73961 298372 73989
rect 298400 73961 298434 73989
rect 298462 73961 298510 73989
rect 298200 65175 298510 73961
rect 298200 65147 298248 65175
rect 298276 65147 298310 65175
rect 298338 65147 298372 65175
rect 298400 65147 298434 65175
rect 298462 65147 298510 65175
rect 298200 65113 298510 65147
rect 298200 65085 298248 65113
rect 298276 65085 298310 65113
rect 298338 65085 298372 65113
rect 298400 65085 298434 65113
rect 298462 65085 298510 65113
rect 298200 65051 298510 65085
rect 298200 65023 298248 65051
rect 298276 65023 298310 65051
rect 298338 65023 298372 65051
rect 298400 65023 298434 65051
rect 298462 65023 298510 65051
rect 298200 64989 298510 65023
rect 298200 64961 298248 64989
rect 298276 64961 298310 64989
rect 298338 64961 298372 64989
rect 298400 64961 298434 64989
rect 298462 64961 298510 64989
rect 298200 56175 298510 64961
rect 298200 56147 298248 56175
rect 298276 56147 298310 56175
rect 298338 56147 298372 56175
rect 298400 56147 298434 56175
rect 298462 56147 298510 56175
rect 298200 56113 298510 56147
rect 298200 56085 298248 56113
rect 298276 56085 298310 56113
rect 298338 56085 298372 56113
rect 298400 56085 298434 56113
rect 298462 56085 298510 56113
rect 298200 56051 298510 56085
rect 298200 56023 298248 56051
rect 298276 56023 298310 56051
rect 298338 56023 298372 56051
rect 298400 56023 298434 56051
rect 298462 56023 298510 56051
rect 298200 55989 298510 56023
rect 298200 55961 298248 55989
rect 298276 55961 298310 55989
rect 298338 55961 298372 55989
rect 298400 55961 298434 55989
rect 298462 55961 298510 55989
rect 298200 47175 298510 55961
rect 298200 47147 298248 47175
rect 298276 47147 298310 47175
rect 298338 47147 298372 47175
rect 298400 47147 298434 47175
rect 298462 47147 298510 47175
rect 298200 47113 298510 47147
rect 298200 47085 298248 47113
rect 298276 47085 298310 47113
rect 298338 47085 298372 47113
rect 298400 47085 298434 47113
rect 298462 47085 298510 47113
rect 298200 47051 298510 47085
rect 298200 47023 298248 47051
rect 298276 47023 298310 47051
rect 298338 47023 298372 47051
rect 298400 47023 298434 47051
rect 298462 47023 298510 47051
rect 298200 46989 298510 47023
rect 298200 46961 298248 46989
rect 298276 46961 298310 46989
rect 298338 46961 298372 46989
rect 298400 46961 298434 46989
rect 298462 46961 298510 46989
rect 298200 38175 298510 46961
rect 298200 38147 298248 38175
rect 298276 38147 298310 38175
rect 298338 38147 298372 38175
rect 298400 38147 298434 38175
rect 298462 38147 298510 38175
rect 298200 38113 298510 38147
rect 298200 38085 298248 38113
rect 298276 38085 298310 38113
rect 298338 38085 298372 38113
rect 298400 38085 298434 38113
rect 298462 38085 298510 38113
rect 298200 38051 298510 38085
rect 298200 38023 298248 38051
rect 298276 38023 298310 38051
rect 298338 38023 298372 38051
rect 298400 38023 298434 38051
rect 298462 38023 298510 38051
rect 298200 37989 298510 38023
rect 298200 37961 298248 37989
rect 298276 37961 298310 37989
rect 298338 37961 298372 37989
rect 298400 37961 298434 37989
rect 298462 37961 298510 37989
rect 298200 29175 298510 37961
rect 298200 29147 298248 29175
rect 298276 29147 298310 29175
rect 298338 29147 298372 29175
rect 298400 29147 298434 29175
rect 298462 29147 298510 29175
rect 298200 29113 298510 29147
rect 298200 29085 298248 29113
rect 298276 29085 298310 29113
rect 298338 29085 298372 29113
rect 298400 29085 298434 29113
rect 298462 29085 298510 29113
rect 298200 29051 298510 29085
rect 298200 29023 298248 29051
rect 298276 29023 298310 29051
rect 298338 29023 298372 29051
rect 298400 29023 298434 29051
rect 298462 29023 298510 29051
rect 298200 28989 298510 29023
rect 298200 28961 298248 28989
rect 298276 28961 298310 28989
rect 298338 28961 298372 28989
rect 298400 28961 298434 28989
rect 298462 28961 298510 28989
rect 298200 20175 298510 28961
rect 298200 20147 298248 20175
rect 298276 20147 298310 20175
rect 298338 20147 298372 20175
rect 298400 20147 298434 20175
rect 298462 20147 298510 20175
rect 298200 20113 298510 20147
rect 298200 20085 298248 20113
rect 298276 20085 298310 20113
rect 298338 20085 298372 20113
rect 298400 20085 298434 20113
rect 298462 20085 298510 20113
rect 298200 20051 298510 20085
rect 298200 20023 298248 20051
rect 298276 20023 298310 20051
rect 298338 20023 298372 20051
rect 298400 20023 298434 20051
rect 298462 20023 298510 20051
rect 298200 19989 298510 20023
rect 298200 19961 298248 19989
rect 298276 19961 298310 19989
rect 298338 19961 298372 19989
rect 298400 19961 298434 19989
rect 298462 19961 298510 19989
rect 298200 11175 298510 19961
rect 298200 11147 298248 11175
rect 298276 11147 298310 11175
rect 298338 11147 298372 11175
rect 298400 11147 298434 11175
rect 298462 11147 298510 11175
rect 298200 11113 298510 11147
rect 298200 11085 298248 11113
rect 298276 11085 298310 11113
rect 298338 11085 298372 11113
rect 298400 11085 298434 11113
rect 298462 11085 298510 11113
rect 298200 11051 298510 11085
rect 298200 11023 298248 11051
rect 298276 11023 298310 11051
rect 298338 11023 298372 11051
rect 298400 11023 298434 11051
rect 298462 11023 298510 11051
rect 298200 10989 298510 11023
rect 298200 10961 298248 10989
rect 298276 10961 298310 10989
rect 298338 10961 298372 10989
rect 298400 10961 298434 10989
rect 298462 10961 298510 10989
rect 298200 2175 298510 10961
rect 298200 2147 298248 2175
rect 298276 2147 298310 2175
rect 298338 2147 298372 2175
rect 298400 2147 298434 2175
rect 298462 2147 298510 2175
rect 298200 2113 298510 2147
rect 298200 2085 298248 2113
rect 298276 2085 298310 2113
rect 298338 2085 298372 2113
rect 298400 2085 298434 2113
rect 298462 2085 298510 2113
rect 298200 2051 298510 2085
rect 298200 2023 298248 2051
rect 298276 2023 298310 2051
rect 298338 2023 298372 2051
rect 298400 2023 298434 2051
rect 298462 2023 298510 2051
rect 298200 1989 298510 2023
rect 298200 1961 298248 1989
rect 298276 1961 298310 1989
rect 298338 1961 298372 1989
rect 298400 1961 298434 1989
rect 298462 1961 298510 1989
rect 298200 -80 298510 1961
rect 298200 -108 298248 -80
rect 298276 -108 298310 -80
rect 298338 -108 298372 -80
rect 298400 -108 298434 -80
rect 298462 -108 298510 -80
rect 298200 -142 298510 -108
rect 298200 -170 298248 -142
rect 298276 -170 298310 -142
rect 298338 -170 298372 -142
rect 298400 -170 298434 -142
rect 298462 -170 298510 -142
rect 298200 -204 298510 -170
rect 298200 -232 298248 -204
rect 298276 -232 298310 -204
rect 298338 -232 298372 -204
rect 298400 -232 298434 -204
rect 298462 -232 298510 -204
rect 298200 -266 298510 -232
rect 298200 -294 298248 -266
rect 298276 -294 298310 -266
rect 298338 -294 298372 -266
rect 298400 -294 298434 -266
rect 298462 -294 298510 -266
rect 298200 -342 298510 -294
rect 298680 293175 298990 298872
rect 298680 293147 298728 293175
rect 298756 293147 298790 293175
rect 298818 293147 298852 293175
rect 298880 293147 298914 293175
rect 298942 293147 298990 293175
rect 298680 293113 298990 293147
rect 298680 293085 298728 293113
rect 298756 293085 298790 293113
rect 298818 293085 298852 293113
rect 298880 293085 298914 293113
rect 298942 293085 298990 293113
rect 298680 293051 298990 293085
rect 298680 293023 298728 293051
rect 298756 293023 298790 293051
rect 298818 293023 298852 293051
rect 298880 293023 298914 293051
rect 298942 293023 298990 293051
rect 298680 292989 298990 293023
rect 298680 292961 298728 292989
rect 298756 292961 298790 292989
rect 298818 292961 298852 292989
rect 298880 292961 298914 292989
rect 298942 292961 298990 292989
rect 298680 284175 298990 292961
rect 298680 284147 298728 284175
rect 298756 284147 298790 284175
rect 298818 284147 298852 284175
rect 298880 284147 298914 284175
rect 298942 284147 298990 284175
rect 298680 284113 298990 284147
rect 298680 284085 298728 284113
rect 298756 284085 298790 284113
rect 298818 284085 298852 284113
rect 298880 284085 298914 284113
rect 298942 284085 298990 284113
rect 298680 284051 298990 284085
rect 298680 284023 298728 284051
rect 298756 284023 298790 284051
rect 298818 284023 298852 284051
rect 298880 284023 298914 284051
rect 298942 284023 298990 284051
rect 298680 283989 298990 284023
rect 298680 283961 298728 283989
rect 298756 283961 298790 283989
rect 298818 283961 298852 283989
rect 298880 283961 298914 283989
rect 298942 283961 298990 283989
rect 298680 275175 298990 283961
rect 298680 275147 298728 275175
rect 298756 275147 298790 275175
rect 298818 275147 298852 275175
rect 298880 275147 298914 275175
rect 298942 275147 298990 275175
rect 298680 275113 298990 275147
rect 298680 275085 298728 275113
rect 298756 275085 298790 275113
rect 298818 275085 298852 275113
rect 298880 275085 298914 275113
rect 298942 275085 298990 275113
rect 298680 275051 298990 275085
rect 298680 275023 298728 275051
rect 298756 275023 298790 275051
rect 298818 275023 298852 275051
rect 298880 275023 298914 275051
rect 298942 275023 298990 275051
rect 298680 274989 298990 275023
rect 298680 274961 298728 274989
rect 298756 274961 298790 274989
rect 298818 274961 298852 274989
rect 298880 274961 298914 274989
rect 298942 274961 298990 274989
rect 298680 266175 298990 274961
rect 298680 266147 298728 266175
rect 298756 266147 298790 266175
rect 298818 266147 298852 266175
rect 298880 266147 298914 266175
rect 298942 266147 298990 266175
rect 298680 266113 298990 266147
rect 298680 266085 298728 266113
rect 298756 266085 298790 266113
rect 298818 266085 298852 266113
rect 298880 266085 298914 266113
rect 298942 266085 298990 266113
rect 298680 266051 298990 266085
rect 298680 266023 298728 266051
rect 298756 266023 298790 266051
rect 298818 266023 298852 266051
rect 298880 266023 298914 266051
rect 298942 266023 298990 266051
rect 298680 265989 298990 266023
rect 298680 265961 298728 265989
rect 298756 265961 298790 265989
rect 298818 265961 298852 265989
rect 298880 265961 298914 265989
rect 298942 265961 298990 265989
rect 298680 257175 298990 265961
rect 298680 257147 298728 257175
rect 298756 257147 298790 257175
rect 298818 257147 298852 257175
rect 298880 257147 298914 257175
rect 298942 257147 298990 257175
rect 298680 257113 298990 257147
rect 298680 257085 298728 257113
rect 298756 257085 298790 257113
rect 298818 257085 298852 257113
rect 298880 257085 298914 257113
rect 298942 257085 298990 257113
rect 298680 257051 298990 257085
rect 298680 257023 298728 257051
rect 298756 257023 298790 257051
rect 298818 257023 298852 257051
rect 298880 257023 298914 257051
rect 298942 257023 298990 257051
rect 298680 256989 298990 257023
rect 298680 256961 298728 256989
rect 298756 256961 298790 256989
rect 298818 256961 298852 256989
rect 298880 256961 298914 256989
rect 298942 256961 298990 256989
rect 298680 248175 298990 256961
rect 298680 248147 298728 248175
rect 298756 248147 298790 248175
rect 298818 248147 298852 248175
rect 298880 248147 298914 248175
rect 298942 248147 298990 248175
rect 298680 248113 298990 248147
rect 298680 248085 298728 248113
rect 298756 248085 298790 248113
rect 298818 248085 298852 248113
rect 298880 248085 298914 248113
rect 298942 248085 298990 248113
rect 298680 248051 298990 248085
rect 298680 248023 298728 248051
rect 298756 248023 298790 248051
rect 298818 248023 298852 248051
rect 298880 248023 298914 248051
rect 298942 248023 298990 248051
rect 298680 247989 298990 248023
rect 298680 247961 298728 247989
rect 298756 247961 298790 247989
rect 298818 247961 298852 247989
rect 298880 247961 298914 247989
rect 298942 247961 298990 247989
rect 298680 239175 298990 247961
rect 298680 239147 298728 239175
rect 298756 239147 298790 239175
rect 298818 239147 298852 239175
rect 298880 239147 298914 239175
rect 298942 239147 298990 239175
rect 298680 239113 298990 239147
rect 298680 239085 298728 239113
rect 298756 239085 298790 239113
rect 298818 239085 298852 239113
rect 298880 239085 298914 239113
rect 298942 239085 298990 239113
rect 298680 239051 298990 239085
rect 298680 239023 298728 239051
rect 298756 239023 298790 239051
rect 298818 239023 298852 239051
rect 298880 239023 298914 239051
rect 298942 239023 298990 239051
rect 298680 238989 298990 239023
rect 298680 238961 298728 238989
rect 298756 238961 298790 238989
rect 298818 238961 298852 238989
rect 298880 238961 298914 238989
rect 298942 238961 298990 238989
rect 298680 230175 298990 238961
rect 298680 230147 298728 230175
rect 298756 230147 298790 230175
rect 298818 230147 298852 230175
rect 298880 230147 298914 230175
rect 298942 230147 298990 230175
rect 298680 230113 298990 230147
rect 298680 230085 298728 230113
rect 298756 230085 298790 230113
rect 298818 230085 298852 230113
rect 298880 230085 298914 230113
rect 298942 230085 298990 230113
rect 298680 230051 298990 230085
rect 298680 230023 298728 230051
rect 298756 230023 298790 230051
rect 298818 230023 298852 230051
rect 298880 230023 298914 230051
rect 298942 230023 298990 230051
rect 298680 229989 298990 230023
rect 298680 229961 298728 229989
rect 298756 229961 298790 229989
rect 298818 229961 298852 229989
rect 298880 229961 298914 229989
rect 298942 229961 298990 229989
rect 298680 221175 298990 229961
rect 298680 221147 298728 221175
rect 298756 221147 298790 221175
rect 298818 221147 298852 221175
rect 298880 221147 298914 221175
rect 298942 221147 298990 221175
rect 298680 221113 298990 221147
rect 298680 221085 298728 221113
rect 298756 221085 298790 221113
rect 298818 221085 298852 221113
rect 298880 221085 298914 221113
rect 298942 221085 298990 221113
rect 298680 221051 298990 221085
rect 298680 221023 298728 221051
rect 298756 221023 298790 221051
rect 298818 221023 298852 221051
rect 298880 221023 298914 221051
rect 298942 221023 298990 221051
rect 298680 220989 298990 221023
rect 298680 220961 298728 220989
rect 298756 220961 298790 220989
rect 298818 220961 298852 220989
rect 298880 220961 298914 220989
rect 298942 220961 298990 220989
rect 298680 212175 298990 220961
rect 298680 212147 298728 212175
rect 298756 212147 298790 212175
rect 298818 212147 298852 212175
rect 298880 212147 298914 212175
rect 298942 212147 298990 212175
rect 298680 212113 298990 212147
rect 298680 212085 298728 212113
rect 298756 212085 298790 212113
rect 298818 212085 298852 212113
rect 298880 212085 298914 212113
rect 298942 212085 298990 212113
rect 298680 212051 298990 212085
rect 298680 212023 298728 212051
rect 298756 212023 298790 212051
rect 298818 212023 298852 212051
rect 298880 212023 298914 212051
rect 298942 212023 298990 212051
rect 298680 211989 298990 212023
rect 298680 211961 298728 211989
rect 298756 211961 298790 211989
rect 298818 211961 298852 211989
rect 298880 211961 298914 211989
rect 298942 211961 298990 211989
rect 298680 203175 298990 211961
rect 298680 203147 298728 203175
rect 298756 203147 298790 203175
rect 298818 203147 298852 203175
rect 298880 203147 298914 203175
rect 298942 203147 298990 203175
rect 298680 203113 298990 203147
rect 298680 203085 298728 203113
rect 298756 203085 298790 203113
rect 298818 203085 298852 203113
rect 298880 203085 298914 203113
rect 298942 203085 298990 203113
rect 298680 203051 298990 203085
rect 298680 203023 298728 203051
rect 298756 203023 298790 203051
rect 298818 203023 298852 203051
rect 298880 203023 298914 203051
rect 298942 203023 298990 203051
rect 298680 202989 298990 203023
rect 298680 202961 298728 202989
rect 298756 202961 298790 202989
rect 298818 202961 298852 202989
rect 298880 202961 298914 202989
rect 298942 202961 298990 202989
rect 298680 194175 298990 202961
rect 298680 194147 298728 194175
rect 298756 194147 298790 194175
rect 298818 194147 298852 194175
rect 298880 194147 298914 194175
rect 298942 194147 298990 194175
rect 298680 194113 298990 194147
rect 298680 194085 298728 194113
rect 298756 194085 298790 194113
rect 298818 194085 298852 194113
rect 298880 194085 298914 194113
rect 298942 194085 298990 194113
rect 298680 194051 298990 194085
rect 298680 194023 298728 194051
rect 298756 194023 298790 194051
rect 298818 194023 298852 194051
rect 298880 194023 298914 194051
rect 298942 194023 298990 194051
rect 298680 193989 298990 194023
rect 298680 193961 298728 193989
rect 298756 193961 298790 193989
rect 298818 193961 298852 193989
rect 298880 193961 298914 193989
rect 298942 193961 298990 193989
rect 298680 185175 298990 193961
rect 298680 185147 298728 185175
rect 298756 185147 298790 185175
rect 298818 185147 298852 185175
rect 298880 185147 298914 185175
rect 298942 185147 298990 185175
rect 298680 185113 298990 185147
rect 298680 185085 298728 185113
rect 298756 185085 298790 185113
rect 298818 185085 298852 185113
rect 298880 185085 298914 185113
rect 298942 185085 298990 185113
rect 298680 185051 298990 185085
rect 298680 185023 298728 185051
rect 298756 185023 298790 185051
rect 298818 185023 298852 185051
rect 298880 185023 298914 185051
rect 298942 185023 298990 185051
rect 298680 184989 298990 185023
rect 298680 184961 298728 184989
rect 298756 184961 298790 184989
rect 298818 184961 298852 184989
rect 298880 184961 298914 184989
rect 298942 184961 298990 184989
rect 298680 176175 298990 184961
rect 298680 176147 298728 176175
rect 298756 176147 298790 176175
rect 298818 176147 298852 176175
rect 298880 176147 298914 176175
rect 298942 176147 298990 176175
rect 298680 176113 298990 176147
rect 298680 176085 298728 176113
rect 298756 176085 298790 176113
rect 298818 176085 298852 176113
rect 298880 176085 298914 176113
rect 298942 176085 298990 176113
rect 298680 176051 298990 176085
rect 298680 176023 298728 176051
rect 298756 176023 298790 176051
rect 298818 176023 298852 176051
rect 298880 176023 298914 176051
rect 298942 176023 298990 176051
rect 298680 175989 298990 176023
rect 298680 175961 298728 175989
rect 298756 175961 298790 175989
rect 298818 175961 298852 175989
rect 298880 175961 298914 175989
rect 298942 175961 298990 175989
rect 298680 167175 298990 175961
rect 298680 167147 298728 167175
rect 298756 167147 298790 167175
rect 298818 167147 298852 167175
rect 298880 167147 298914 167175
rect 298942 167147 298990 167175
rect 298680 167113 298990 167147
rect 298680 167085 298728 167113
rect 298756 167085 298790 167113
rect 298818 167085 298852 167113
rect 298880 167085 298914 167113
rect 298942 167085 298990 167113
rect 298680 167051 298990 167085
rect 298680 167023 298728 167051
rect 298756 167023 298790 167051
rect 298818 167023 298852 167051
rect 298880 167023 298914 167051
rect 298942 167023 298990 167051
rect 298680 166989 298990 167023
rect 298680 166961 298728 166989
rect 298756 166961 298790 166989
rect 298818 166961 298852 166989
rect 298880 166961 298914 166989
rect 298942 166961 298990 166989
rect 298680 158175 298990 166961
rect 298680 158147 298728 158175
rect 298756 158147 298790 158175
rect 298818 158147 298852 158175
rect 298880 158147 298914 158175
rect 298942 158147 298990 158175
rect 298680 158113 298990 158147
rect 298680 158085 298728 158113
rect 298756 158085 298790 158113
rect 298818 158085 298852 158113
rect 298880 158085 298914 158113
rect 298942 158085 298990 158113
rect 298680 158051 298990 158085
rect 298680 158023 298728 158051
rect 298756 158023 298790 158051
rect 298818 158023 298852 158051
rect 298880 158023 298914 158051
rect 298942 158023 298990 158051
rect 298680 157989 298990 158023
rect 298680 157961 298728 157989
rect 298756 157961 298790 157989
rect 298818 157961 298852 157989
rect 298880 157961 298914 157989
rect 298942 157961 298990 157989
rect 298680 149175 298990 157961
rect 298680 149147 298728 149175
rect 298756 149147 298790 149175
rect 298818 149147 298852 149175
rect 298880 149147 298914 149175
rect 298942 149147 298990 149175
rect 298680 149113 298990 149147
rect 298680 149085 298728 149113
rect 298756 149085 298790 149113
rect 298818 149085 298852 149113
rect 298880 149085 298914 149113
rect 298942 149085 298990 149113
rect 298680 149051 298990 149085
rect 298680 149023 298728 149051
rect 298756 149023 298790 149051
rect 298818 149023 298852 149051
rect 298880 149023 298914 149051
rect 298942 149023 298990 149051
rect 298680 148989 298990 149023
rect 298680 148961 298728 148989
rect 298756 148961 298790 148989
rect 298818 148961 298852 148989
rect 298880 148961 298914 148989
rect 298942 148961 298990 148989
rect 298680 140175 298990 148961
rect 298680 140147 298728 140175
rect 298756 140147 298790 140175
rect 298818 140147 298852 140175
rect 298880 140147 298914 140175
rect 298942 140147 298990 140175
rect 298680 140113 298990 140147
rect 298680 140085 298728 140113
rect 298756 140085 298790 140113
rect 298818 140085 298852 140113
rect 298880 140085 298914 140113
rect 298942 140085 298990 140113
rect 298680 140051 298990 140085
rect 298680 140023 298728 140051
rect 298756 140023 298790 140051
rect 298818 140023 298852 140051
rect 298880 140023 298914 140051
rect 298942 140023 298990 140051
rect 298680 139989 298990 140023
rect 298680 139961 298728 139989
rect 298756 139961 298790 139989
rect 298818 139961 298852 139989
rect 298880 139961 298914 139989
rect 298942 139961 298990 139989
rect 298680 131175 298990 139961
rect 298680 131147 298728 131175
rect 298756 131147 298790 131175
rect 298818 131147 298852 131175
rect 298880 131147 298914 131175
rect 298942 131147 298990 131175
rect 298680 131113 298990 131147
rect 298680 131085 298728 131113
rect 298756 131085 298790 131113
rect 298818 131085 298852 131113
rect 298880 131085 298914 131113
rect 298942 131085 298990 131113
rect 298680 131051 298990 131085
rect 298680 131023 298728 131051
rect 298756 131023 298790 131051
rect 298818 131023 298852 131051
rect 298880 131023 298914 131051
rect 298942 131023 298990 131051
rect 298680 130989 298990 131023
rect 298680 130961 298728 130989
rect 298756 130961 298790 130989
rect 298818 130961 298852 130989
rect 298880 130961 298914 130989
rect 298942 130961 298990 130989
rect 298680 122175 298990 130961
rect 298680 122147 298728 122175
rect 298756 122147 298790 122175
rect 298818 122147 298852 122175
rect 298880 122147 298914 122175
rect 298942 122147 298990 122175
rect 298680 122113 298990 122147
rect 298680 122085 298728 122113
rect 298756 122085 298790 122113
rect 298818 122085 298852 122113
rect 298880 122085 298914 122113
rect 298942 122085 298990 122113
rect 298680 122051 298990 122085
rect 298680 122023 298728 122051
rect 298756 122023 298790 122051
rect 298818 122023 298852 122051
rect 298880 122023 298914 122051
rect 298942 122023 298990 122051
rect 298680 121989 298990 122023
rect 298680 121961 298728 121989
rect 298756 121961 298790 121989
rect 298818 121961 298852 121989
rect 298880 121961 298914 121989
rect 298942 121961 298990 121989
rect 298680 113175 298990 121961
rect 298680 113147 298728 113175
rect 298756 113147 298790 113175
rect 298818 113147 298852 113175
rect 298880 113147 298914 113175
rect 298942 113147 298990 113175
rect 298680 113113 298990 113147
rect 298680 113085 298728 113113
rect 298756 113085 298790 113113
rect 298818 113085 298852 113113
rect 298880 113085 298914 113113
rect 298942 113085 298990 113113
rect 298680 113051 298990 113085
rect 298680 113023 298728 113051
rect 298756 113023 298790 113051
rect 298818 113023 298852 113051
rect 298880 113023 298914 113051
rect 298942 113023 298990 113051
rect 298680 112989 298990 113023
rect 298680 112961 298728 112989
rect 298756 112961 298790 112989
rect 298818 112961 298852 112989
rect 298880 112961 298914 112989
rect 298942 112961 298990 112989
rect 298680 104175 298990 112961
rect 298680 104147 298728 104175
rect 298756 104147 298790 104175
rect 298818 104147 298852 104175
rect 298880 104147 298914 104175
rect 298942 104147 298990 104175
rect 298680 104113 298990 104147
rect 298680 104085 298728 104113
rect 298756 104085 298790 104113
rect 298818 104085 298852 104113
rect 298880 104085 298914 104113
rect 298942 104085 298990 104113
rect 298680 104051 298990 104085
rect 298680 104023 298728 104051
rect 298756 104023 298790 104051
rect 298818 104023 298852 104051
rect 298880 104023 298914 104051
rect 298942 104023 298990 104051
rect 298680 103989 298990 104023
rect 298680 103961 298728 103989
rect 298756 103961 298790 103989
rect 298818 103961 298852 103989
rect 298880 103961 298914 103989
rect 298942 103961 298990 103989
rect 298680 95175 298990 103961
rect 298680 95147 298728 95175
rect 298756 95147 298790 95175
rect 298818 95147 298852 95175
rect 298880 95147 298914 95175
rect 298942 95147 298990 95175
rect 298680 95113 298990 95147
rect 298680 95085 298728 95113
rect 298756 95085 298790 95113
rect 298818 95085 298852 95113
rect 298880 95085 298914 95113
rect 298942 95085 298990 95113
rect 298680 95051 298990 95085
rect 298680 95023 298728 95051
rect 298756 95023 298790 95051
rect 298818 95023 298852 95051
rect 298880 95023 298914 95051
rect 298942 95023 298990 95051
rect 298680 94989 298990 95023
rect 298680 94961 298728 94989
rect 298756 94961 298790 94989
rect 298818 94961 298852 94989
rect 298880 94961 298914 94989
rect 298942 94961 298990 94989
rect 298680 86175 298990 94961
rect 298680 86147 298728 86175
rect 298756 86147 298790 86175
rect 298818 86147 298852 86175
rect 298880 86147 298914 86175
rect 298942 86147 298990 86175
rect 298680 86113 298990 86147
rect 298680 86085 298728 86113
rect 298756 86085 298790 86113
rect 298818 86085 298852 86113
rect 298880 86085 298914 86113
rect 298942 86085 298990 86113
rect 298680 86051 298990 86085
rect 298680 86023 298728 86051
rect 298756 86023 298790 86051
rect 298818 86023 298852 86051
rect 298880 86023 298914 86051
rect 298942 86023 298990 86051
rect 298680 85989 298990 86023
rect 298680 85961 298728 85989
rect 298756 85961 298790 85989
rect 298818 85961 298852 85989
rect 298880 85961 298914 85989
rect 298942 85961 298990 85989
rect 298680 77175 298990 85961
rect 298680 77147 298728 77175
rect 298756 77147 298790 77175
rect 298818 77147 298852 77175
rect 298880 77147 298914 77175
rect 298942 77147 298990 77175
rect 298680 77113 298990 77147
rect 298680 77085 298728 77113
rect 298756 77085 298790 77113
rect 298818 77085 298852 77113
rect 298880 77085 298914 77113
rect 298942 77085 298990 77113
rect 298680 77051 298990 77085
rect 298680 77023 298728 77051
rect 298756 77023 298790 77051
rect 298818 77023 298852 77051
rect 298880 77023 298914 77051
rect 298942 77023 298990 77051
rect 298680 76989 298990 77023
rect 298680 76961 298728 76989
rect 298756 76961 298790 76989
rect 298818 76961 298852 76989
rect 298880 76961 298914 76989
rect 298942 76961 298990 76989
rect 298680 68175 298990 76961
rect 298680 68147 298728 68175
rect 298756 68147 298790 68175
rect 298818 68147 298852 68175
rect 298880 68147 298914 68175
rect 298942 68147 298990 68175
rect 298680 68113 298990 68147
rect 298680 68085 298728 68113
rect 298756 68085 298790 68113
rect 298818 68085 298852 68113
rect 298880 68085 298914 68113
rect 298942 68085 298990 68113
rect 298680 68051 298990 68085
rect 298680 68023 298728 68051
rect 298756 68023 298790 68051
rect 298818 68023 298852 68051
rect 298880 68023 298914 68051
rect 298942 68023 298990 68051
rect 298680 67989 298990 68023
rect 298680 67961 298728 67989
rect 298756 67961 298790 67989
rect 298818 67961 298852 67989
rect 298880 67961 298914 67989
rect 298942 67961 298990 67989
rect 298680 59175 298990 67961
rect 298680 59147 298728 59175
rect 298756 59147 298790 59175
rect 298818 59147 298852 59175
rect 298880 59147 298914 59175
rect 298942 59147 298990 59175
rect 298680 59113 298990 59147
rect 298680 59085 298728 59113
rect 298756 59085 298790 59113
rect 298818 59085 298852 59113
rect 298880 59085 298914 59113
rect 298942 59085 298990 59113
rect 298680 59051 298990 59085
rect 298680 59023 298728 59051
rect 298756 59023 298790 59051
rect 298818 59023 298852 59051
rect 298880 59023 298914 59051
rect 298942 59023 298990 59051
rect 298680 58989 298990 59023
rect 298680 58961 298728 58989
rect 298756 58961 298790 58989
rect 298818 58961 298852 58989
rect 298880 58961 298914 58989
rect 298942 58961 298990 58989
rect 298680 50175 298990 58961
rect 298680 50147 298728 50175
rect 298756 50147 298790 50175
rect 298818 50147 298852 50175
rect 298880 50147 298914 50175
rect 298942 50147 298990 50175
rect 298680 50113 298990 50147
rect 298680 50085 298728 50113
rect 298756 50085 298790 50113
rect 298818 50085 298852 50113
rect 298880 50085 298914 50113
rect 298942 50085 298990 50113
rect 298680 50051 298990 50085
rect 298680 50023 298728 50051
rect 298756 50023 298790 50051
rect 298818 50023 298852 50051
rect 298880 50023 298914 50051
rect 298942 50023 298990 50051
rect 298680 49989 298990 50023
rect 298680 49961 298728 49989
rect 298756 49961 298790 49989
rect 298818 49961 298852 49989
rect 298880 49961 298914 49989
rect 298942 49961 298990 49989
rect 298680 41175 298990 49961
rect 298680 41147 298728 41175
rect 298756 41147 298790 41175
rect 298818 41147 298852 41175
rect 298880 41147 298914 41175
rect 298942 41147 298990 41175
rect 298680 41113 298990 41147
rect 298680 41085 298728 41113
rect 298756 41085 298790 41113
rect 298818 41085 298852 41113
rect 298880 41085 298914 41113
rect 298942 41085 298990 41113
rect 298680 41051 298990 41085
rect 298680 41023 298728 41051
rect 298756 41023 298790 41051
rect 298818 41023 298852 41051
rect 298880 41023 298914 41051
rect 298942 41023 298990 41051
rect 298680 40989 298990 41023
rect 298680 40961 298728 40989
rect 298756 40961 298790 40989
rect 298818 40961 298852 40989
rect 298880 40961 298914 40989
rect 298942 40961 298990 40989
rect 298680 32175 298990 40961
rect 298680 32147 298728 32175
rect 298756 32147 298790 32175
rect 298818 32147 298852 32175
rect 298880 32147 298914 32175
rect 298942 32147 298990 32175
rect 298680 32113 298990 32147
rect 298680 32085 298728 32113
rect 298756 32085 298790 32113
rect 298818 32085 298852 32113
rect 298880 32085 298914 32113
rect 298942 32085 298990 32113
rect 298680 32051 298990 32085
rect 298680 32023 298728 32051
rect 298756 32023 298790 32051
rect 298818 32023 298852 32051
rect 298880 32023 298914 32051
rect 298942 32023 298990 32051
rect 298680 31989 298990 32023
rect 298680 31961 298728 31989
rect 298756 31961 298790 31989
rect 298818 31961 298852 31989
rect 298880 31961 298914 31989
rect 298942 31961 298990 31989
rect 298680 23175 298990 31961
rect 298680 23147 298728 23175
rect 298756 23147 298790 23175
rect 298818 23147 298852 23175
rect 298880 23147 298914 23175
rect 298942 23147 298990 23175
rect 298680 23113 298990 23147
rect 298680 23085 298728 23113
rect 298756 23085 298790 23113
rect 298818 23085 298852 23113
rect 298880 23085 298914 23113
rect 298942 23085 298990 23113
rect 298680 23051 298990 23085
rect 298680 23023 298728 23051
rect 298756 23023 298790 23051
rect 298818 23023 298852 23051
rect 298880 23023 298914 23051
rect 298942 23023 298990 23051
rect 298680 22989 298990 23023
rect 298680 22961 298728 22989
rect 298756 22961 298790 22989
rect 298818 22961 298852 22989
rect 298880 22961 298914 22989
rect 298942 22961 298990 22989
rect 298680 14175 298990 22961
rect 298680 14147 298728 14175
rect 298756 14147 298790 14175
rect 298818 14147 298852 14175
rect 298880 14147 298914 14175
rect 298942 14147 298990 14175
rect 298680 14113 298990 14147
rect 298680 14085 298728 14113
rect 298756 14085 298790 14113
rect 298818 14085 298852 14113
rect 298880 14085 298914 14113
rect 298942 14085 298990 14113
rect 298680 14051 298990 14085
rect 298680 14023 298728 14051
rect 298756 14023 298790 14051
rect 298818 14023 298852 14051
rect 298880 14023 298914 14051
rect 298942 14023 298990 14051
rect 298680 13989 298990 14023
rect 298680 13961 298728 13989
rect 298756 13961 298790 13989
rect 298818 13961 298852 13989
rect 298880 13961 298914 13989
rect 298942 13961 298990 13989
rect 298680 5175 298990 13961
rect 298680 5147 298728 5175
rect 298756 5147 298790 5175
rect 298818 5147 298852 5175
rect 298880 5147 298914 5175
rect 298942 5147 298990 5175
rect 298680 5113 298990 5147
rect 298680 5085 298728 5113
rect 298756 5085 298790 5113
rect 298818 5085 298852 5113
rect 298880 5085 298914 5113
rect 298942 5085 298990 5113
rect 298680 5051 298990 5085
rect 298680 5023 298728 5051
rect 298756 5023 298790 5051
rect 298818 5023 298852 5051
rect 298880 5023 298914 5051
rect 298942 5023 298990 5051
rect 298680 4989 298990 5023
rect 298680 4961 298728 4989
rect 298756 4961 298790 4989
rect 298818 4961 298852 4989
rect 298880 4961 298914 4989
rect 298942 4961 298990 4989
rect 296409 -588 296457 -560
rect 296485 -588 296519 -560
rect 296547 -588 296581 -560
rect 296609 -588 296643 -560
rect 296671 -588 296719 -560
rect 296409 -622 296719 -588
rect 296409 -650 296457 -622
rect 296485 -650 296519 -622
rect 296547 -650 296581 -622
rect 296609 -650 296643 -622
rect 296671 -650 296719 -622
rect 296409 -684 296719 -650
rect 296409 -712 296457 -684
rect 296485 -712 296519 -684
rect 296547 -712 296581 -684
rect 296609 -712 296643 -684
rect 296671 -712 296719 -684
rect 296409 -746 296719 -712
rect 296409 -774 296457 -746
rect 296485 -774 296519 -746
rect 296547 -774 296581 -746
rect 296609 -774 296643 -746
rect 296671 -774 296719 -746
rect 296409 -822 296719 -774
rect 298680 -560 298990 4961
rect 298680 -588 298728 -560
rect 298756 -588 298790 -560
rect 298818 -588 298852 -560
rect 298880 -588 298914 -560
rect 298942 -588 298990 -560
rect 298680 -622 298990 -588
rect 298680 -650 298728 -622
rect 298756 -650 298790 -622
rect 298818 -650 298852 -622
rect 298880 -650 298914 -622
rect 298942 -650 298990 -622
rect 298680 -684 298990 -650
rect 298680 -712 298728 -684
rect 298756 -712 298790 -684
rect 298818 -712 298852 -684
rect 298880 -712 298914 -684
rect 298942 -712 298990 -684
rect 298680 -746 298990 -712
rect 298680 -774 298728 -746
rect 298756 -774 298790 -746
rect 298818 -774 298852 -746
rect 298880 -774 298914 -746
rect 298942 -774 298990 -746
rect 298680 -822 298990 -774
<< via4 >>
rect -910 299058 -882 299086
rect -848 299058 -820 299086
rect -786 299058 -758 299086
rect -724 299058 -696 299086
rect -910 298996 -882 299024
rect -848 298996 -820 299024
rect -786 298996 -758 299024
rect -724 298996 -696 299024
rect -910 298934 -882 298962
rect -848 298934 -820 298962
rect -786 298934 -758 298962
rect -724 298934 -696 298962
rect -910 298872 -882 298900
rect -848 298872 -820 298900
rect -786 298872 -758 298900
rect -724 298872 -696 298900
rect -910 293147 -882 293175
rect -848 293147 -820 293175
rect -786 293147 -758 293175
rect -724 293147 -696 293175
rect -910 293085 -882 293113
rect -848 293085 -820 293113
rect -786 293085 -758 293113
rect -724 293085 -696 293113
rect -910 293023 -882 293051
rect -848 293023 -820 293051
rect -786 293023 -758 293051
rect -724 293023 -696 293051
rect -910 292961 -882 292989
rect -848 292961 -820 292989
rect -786 292961 -758 292989
rect -724 292961 -696 292989
rect -910 284147 -882 284175
rect -848 284147 -820 284175
rect -786 284147 -758 284175
rect -724 284147 -696 284175
rect -910 284085 -882 284113
rect -848 284085 -820 284113
rect -786 284085 -758 284113
rect -724 284085 -696 284113
rect -910 284023 -882 284051
rect -848 284023 -820 284051
rect -786 284023 -758 284051
rect -724 284023 -696 284051
rect -910 283961 -882 283989
rect -848 283961 -820 283989
rect -786 283961 -758 283989
rect -724 283961 -696 283989
rect -910 275147 -882 275175
rect -848 275147 -820 275175
rect -786 275147 -758 275175
rect -724 275147 -696 275175
rect -910 275085 -882 275113
rect -848 275085 -820 275113
rect -786 275085 -758 275113
rect -724 275085 -696 275113
rect -910 275023 -882 275051
rect -848 275023 -820 275051
rect -786 275023 -758 275051
rect -724 275023 -696 275051
rect -910 274961 -882 274989
rect -848 274961 -820 274989
rect -786 274961 -758 274989
rect -724 274961 -696 274989
rect -910 266147 -882 266175
rect -848 266147 -820 266175
rect -786 266147 -758 266175
rect -724 266147 -696 266175
rect -910 266085 -882 266113
rect -848 266085 -820 266113
rect -786 266085 -758 266113
rect -724 266085 -696 266113
rect -910 266023 -882 266051
rect -848 266023 -820 266051
rect -786 266023 -758 266051
rect -724 266023 -696 266051
rect -910 265961 -882 265989
rect -848 265961 -820 265989
rect -786 265961 -758 265989
rect -724 265961 -696 265989
rect -910 257147 -882 257175
rect -848 257147 -820 257175
rect -786 257147 -758 257175
rect -724 257147 -696 257175
rect -910 257085 -882 257113
rect -848 257085 -820 257113
rect -786 257085 -758 257113
rect -724 257085 -696 257113
rect -910 257023 -882 257051
rect -848 257023 -820 257051
rect -786 257023 -758 257051
rect -724 257023 -696 257051
rect -910 256961 -882 256989
rect -848 256961 -820 256989
rect -786 256961 -758 256989
rect -724 256961 -696 256989
rect -910 248147 -882 248175
rect -848 248147 -820 248175
rect -786 248147 -758 248175
rect -724 248147 -696 248175
rect -910 248085 -882 248113
rect -848 248085 -820 248113
rect -786 248085 -758 248113
rect -724 248085 -696 248113
rect -910 248023 -882 248051
rect -848 248023 -820 248051
rect -786 248023 -758 248051
rect -724 248023 -696 248051
rect -910 247961 -882 247989
rect -848 247961 -820 247989
rect -786 247961 -758 247989
rect -724 247961 -696 247989
rect -910 239147 -882 239175
rect -848 239147 -820 239175
rect -786 239147 -758 239175
rect -724 239147 -696 239175
rect -910 239085 -882 239113
rect -848 239085 -820 239113
rect -786 239085 -758 239113
rect -724 239085 -696 239113
rect -910 239023 -882 239051
rect -848 239023 -820 239051
rect -786 239023 -758 239051
rect -724 239023 -696 239051
rect -910 238961 -882 238989
rect -848 238961 -820 238989
rect -786 238961 -758 238989
rect -724 238961 -696 238989
rect -910 230147 -882 230175
rect -848 230147 -820 230175
rect -786 230147 -758 230175
rect -724 230147 -696 230175
rect -910 230085 -882 230113
rect -848 230085 -820 230113
rect -786 230085 -758 230113
rect -724 230085 -696 230113
rect -910 230023 -882 230051
rect -848 230023 -820 230051
rect -786 230023 -758 230051
rect -724 230023 -696 230051
rect -910 229961 -882 229989
rect -848 229961 -820 229989
rect -786 229961 -758 229989
rect -724 229961 -696 229989
rect -910 221147 -882 221175
rect -848 221147 -820 221175
rect -786 221147 -758 221175
rect -724 221147 -696 221175
rect -910 221085 -882 221113
rect -848 221085 -820 221113
rect -786 221085 -758 221113
rect -724 221085 -696 221113
rect -910 221023 -882 221051
rect -848 221023 -820 221051
rect -786 221023 -758 221051
rect -724 221023 -696 221051
rect -910 220961 -882 220989
rect -848 220961 -820 220989
rect -786 220961 -758 220989
rect -724 220961 -696 220989
rect -910 212147 -882 212175
rect -848 212147 -820 212175
rect -786 212147 -758 212175
rect -724 212147 -696 212175
rect -910 212085 -882 212113
rect -848 212085 -820 212113
rect -786 212085 -758 212113
rect -724 212085 -696 212113
rect -910 212023 -882 212051
rect -848 212023 -820 212051
rect -786 212023 -758 212051
rect -724 212023 -696 212051
rect -910 211961 -882 211989
rect -848 211961 -820 211989
rect -786 211961 -758 211989
rect -724 211961 -696 211989
rect -910 203147 -882 203175
rect -848 203147 -820 203175
rect -786 203147 -758 203175
rect -724 203147 -696 203175
rect -910 203085 -882 203113
rect -848 203085 -820 203113
rect -786 203085 -758 203113
rect -724 203085 -696 203113
rect -910 203023 -882 203051
rect -848 203023 -820 203051
rect -786 203023 -758 203051
rect -724 203023 -696 203051
rect -910 202961 -882 202989
rect -848 202961 -820 202989
rect -786 202961 -758 202989
rect -724 202961 -696 202989
rect -910 194147 -882 194175
rect -848 194147 -820 194175
rect -786 194147 -758 194175
rect -724 194147 -696 194175
rect -910 194085 -882 194113
rect -848 194085 -820 194113
rect -786 194085 -758 194113
rect -724 194085 -696 194113
rect -910 194023 -882 194051
rect -848 194023 -820 194051
rect -786 194023 -758 194051
rect -724 194023 -696 194051
rect -910 193961 -882 193989
rect -848 193961 -820 193989
rect -786 193961 -758 193989
rect -724 193961 -696 193989
rect -910 185147 -882 185175
rect -848 185147 -820 185175
rect -786 185147 -758 185175
rect -724 185147 -696 185175
rect -910 185085 -882 185113
rect -848 185085 -820 185113
rect -786 185085 -758 185113
rect -724 185085 -696 185113
rect -910 185023 -882 185051
rect -848 185023 -820 185051
rect -786 185023 -758 185051
rect -724 185023 -696 185051
rect -910 184961 -882 184989
rect -848 184961 -820 184989
rect -786 184961 -758 184989
rect -724 184961 -696 184989
rect -910 176147 -882 176175
rect -848 176147 -820 176175
rect -786 176147 -758 176175
rect -724 176147 -696 176175
rect -910 176085 -882 176113
rect -848 176085 -820 176113
rect -786 176085 -758 176113
rect -724 176085 -696 176113
rect -910 176023 -882 176051
rect -848 176023 -820 176051
rect -786 176023 -758 176051
rect -724 176023 -696 176051
rect -910 175961 -882 175989
rect -848 175961 -820 175989
rect -786 175961 -758 175989
rect -724 175961 -696 175989
rect -910 167147 -882 167175
rect -848 167147 -820 167175
rect -786 167147 -758 167175
rect -724 167147 -696 167175
rect -910 167085 -882 167113
rect -848 167085 -820 167113
rect -786 167085 -758 167113
rect -724 167085 -696 167113
rect -910 167023 -882 167051
rect -848 167023 -820 167051
rect -786 167023 -758 167051
rect -724 167023 -696 167051
rect -910 166961 -882 166989
rect -848 166961 -820 166989
rect -786 166961 -758 166989
rect -724 166961 -696 166989
rect -910 158147 -882 158175
rect -848 158147 -820 158175
rect -786 158147 -758 158175
rect -724 158147 -696 158175
rect -910 158085 -882 158113
rect -848 158085 -820 158113
rect -786 158085 -758 158113
rect -724 158085 -696 158113
rect -910 158023 -882 158051
rect -848 158023 -820 158051
rect -786 158023 -758 158051
rect -724 158023 -696 158051
rect -910 157961 -882 157989
rect -848 157961 -820 157989
rect -786 157961 -758 157989
rect -724 157961 -696 157989
rect -910 149147 -882 149175
rect -848 149147 -820 149175
rect -786 149147 -758 149175
rect -724 149147 -696 149175
rect -910 149085 -882 149113
rect -848 149085 -820 149113
rect -786 149085 -758 149113
rect -724 149085 -696 149113
rect -910 149023 -882 149051
rect -848 149023 -820 149051
rect -786 149023 -758 149051
rect -724 149023 -696 149051
rect -910 148961 -882 148989
rect -848 148961 -820 148989
rect -786 148961 -758 148989
rect -724 148961 -696 148989
rect -910 140147 -882 140175
rect -848 140147 -820 140175
rect -786 140147 -758 140175
rect -724 140147 -696 140175
rect -910 140085 -882 140113
rect -848 140085 -820 140113
rect -786 140085 -758 140113
rect -724 140085 -696 140113
rect -910 140023 -882 140051
rect -848 140023 -820 140051
rect -786 140023 -758 140051
rect -724 140023 -696 140051
rect -910 139961 -882 139989
rect -848 139961 -820 139989
rect -786 139961 -758 139989
rect -724 139961 -696 139989
rect -910 131147 -882 131175
rect -848 131147 -820 131175
rect -786 131147 -758 131175
rect -724 131147 -696 131175
rect -910 131085 -882 131113
rect -848 131085 -820 131113
rect -786 131085 -758 131113
rect -724 131085 -696 131113
rect -910 131023 -882 131051
rect -848 131023 -820 131051
rect -786 131023 -758 131051
rect -724 131023 -696 131051
rect -910 130961 -882 130989
rect -848 130961 -820 130989
rect -786 130961 -758 130989
rect -724 130961 -696 130989
rect -910 122147 -882 122175
rect -848 122147 -820 122175
rect -786 122147 -758 122175
rect -724 122147 -696 122175
rect -910 122085 -882 122113
rect -848 122085 -820 122113
rect -786 122085 -758 122113
rect -724 122085 -696 122113
rect -910 122023 -882 122051
rect -848 122023 -820 122051
rect -786 122023 -758 122051
rect -724 122023 -696 122051
rect -910 121961 -882 121989
rect -848 121961 -820 121989
rect -786 121961 -758 121989
rect -724 121961 -696 121989
rect -910 113147 -882 113175
rect -848 113147 -820 113175
rect -786 113147 -758 113175
rect -724 113147 -696 113175
rect -910 113085 -882 113113
rect -848 113085 -820 113113
rect -786 113085 -758 113113
rect -724 113085 -696 113113
rect -910 113023 -882 113051
rect -848 113023 -820 113051
rect -786 113023 -758 113051
rect -724 113023 -696 113051
rect -910 112961 -882 112989
rect -848 112961 -820 112989
rect -786 112961 -758 112989
rect -724 112961 -696 112989
rect -910 104147 -882 104175
rect -848 104147 -820 104175
rect -786 104147 -758 104175
rect -724 104147 -696 104175
rect -910 104085 -882 104113
rect -848 104085 -820 104113
rect -786 104085 -758 104113
rect -724 104085 -696 104113
rect -910 104023 -882 104051
rect -848 104023 -820 104051
rect -786 104023 -758 104051
rect -724 104023 -696 104051
rect -910 103961 -882 103989
rect -848 103961 -820 103989
rect -786 103961 -758 103989
rect -724 103961 -696 103989
rect -910 95147 -882 95175
rect -848 95147 -820 95175
rect -786 95147 -758 95175
rect -724 95147 -696 95175
rect -910 95085 -882 95113
rect -848 95085 -820 95113
rect -786 95085 -758 95113
rect -724 95085 -696 95113
rect -910 95023 -882 95051
rect -848 95023 -820 95051
rect -786 95023 -758 95051
rect -724 95023 -696 95051
rect -910 94961 -882 94989
rect -848 94961 -820 94989
rect -786 94961 -758 94989
rect -724 94961 -696 94989
rect -910 86147 -882 86175
rect -848 86147 -820 86175
rect -786 86147 -758 86175
rect -724 86147 -696 86175
rect -910 86085 -882 86113
rect -848 86085 -820 86113
rect -786 86085 -758 86113
rect -724 86085 -696 86113
rect -910 86023 -882 86051
rect -848 86023 -820 86051
rect -786 86023 -758 86051
rect -724 86023 -696 86051
rect -910 85961 -882 85989
rect -848 85961 -820 85989
rect -786 85961 -758 85989
rect -724 85961 -696 85989
rect -910 77147 -882 77175
rect -848 77147 -820 77175
rect -786 77147 -758 77175
rect -724 77147 -696 77175
rect -910 77085 -882 77113
rect -848 77085 -820 77113
rect -786 77085 -758 77113
rect -724 77085 -696 77113
rect -910 77023 -882 77051
rect -848 77023 -820 77051
rect -786 77023 -758 77051
rect -724 77023 -696 77051
rect -910 76961 -882 76989
rect -848 76961 -820 76989
rect -786 76961 -758 76989
rect -724 76961 -696 76989
rect -910 68147 -882 68175
rect -848 68147 -820 68175
rect -786 68147 -758 68175
rect -724 68147 -696 68175
rect -910 68085 -882 68113
rect -848 68085 -820 68113
rect -786 68085 -758 68113
rect -724 68085 -696 68113
rect -910 68023 -882 68051
rect -848 68023 -820 68051
rect -786 68023 -758 68051
rect -724 68023 -696 68051
rect -910 67961 -882 67989
rect -848 67961 -820 67989
rect -786 67961 -758 67989
rect -724 67961 -696 67989
rect -910 59147 -882 59175
rect -848 59147 -820 59175
rect -786 59147 -758 59175
rect -724 59147 -696 59175
rect -910 59085 -882 59113
rect -848 59085 -820 59113
rect -786 59085 -758 59113
rect -724 59085 -696 59113
rect -910 59023 -882 59051
rect -848 59023 -820 59051
rect -786 59023 -758 59051
rect -724 59023 -696 59051
rect -910 58961 -882 58989
rect -848 58961 -820 58989
rect -786 58961 -758 58989
rect -724 58961 -696 58989
rect -910 50147 -882 50175
rect -848 50147 -820 50175
rect -786 50147 -758 50175
rect -724 50147 -696 50175
rect -910 50085 -882 50113
rect -848 50085 -820 50113
rect -786 50085 -758 50113
rect -724 50085 -696 50113
rect -910 50023 -882 50051
rect -848 50023 -820 50051
rect -786 50023 -758 50051
rect -724 50023 -696 50051
rect -910 49961 -882 49989
rect -848 49961 -820 49989
rect -786 49961 -758 49989
rect -724 49961 -696 49989
rect -910 41147 -882 41175
rect -848 41147 -820 41175
rect -786 41147 -758 41175
rect -724 41147 -696 41175
rect -910 41085 -882 41113
rect -848 41085 -820 41113
rect -786 41085 -758 41113
rect -724 41085 -696 41113
rect -910 41023 -882 41051
rect -848 41023 -820 41051
rect -786 41023 -758 41051
rect -724 41023 -696 41051
rect -910 40961 -882 40989
rect -848 40961 -820 40989
rect -786 40961 -758 40989
rect -724 40961 -696 40989
rect -910 32147 -882 32175
rect -848 32147 -820 32175
rect -786 32147 -758 32175
rect -724 32147 -696 32175
rect -910 32085 -882 32113
rect -848 32085 -820 32113
rect -786 32085 -758 32113
rect -724 32085 -696 32113
rect -910 32023 -882 32051
rect -848 32023 -820 32051
rect -786 32023 -758 32051
rect -724 32023 -696 32051
rect -910 31961 -882 31989
rect -848 31961 -820 31989
rect -786 31961 -758 31989
rect -724 31961 -696 31989
rect -910 23147 -882 23175
rect -848 23147 -820 23175
rect -786 23147 -758 23175
rect -724 23147 -696 23175
rect -910 23085 -882 23113
rect -848 23085 -820 23113
rect -786 23085 -758 23113
rect -724 23085 -696 23113
rect -910 23023 -882 23051
rect -848 23023 -820 23051
rect -786 23023 -758 23051
rect -724 23023 -696 23051
rect -910 22961 -882 22989
rect -848 22961 -820 22989
rect -786 22961 -758 22989
rect -724 22961 -696 22989
rect -910 14147 -882 14175
rect -848 14147 -820 14175
rect -786 14147 -758 14175
rect -724 14147 -696 14175
rect -910 14085 -882 14113
rect -848 14085 -820 14113
rect -786 14085 -758 14113
rect -724 14085 -696 14113
rect -910 14023 -882 14051
rect -848 14023 -820 14051
rect -786 14023 -758 14051
rect -724 14023 -696 14051
rect -910 13961 -882 13989
rect -848 13961 -820 13989
rect -786 13961 -758 13989
rect -724 13961 -696 13989
rect -910 5147 -882 5175
rect -848 5147 -820 5175
rect -786 5147 -758 5175
rect -724 5147 -696 5175
rect -910 5085 -882 5113
rect -848 5085 -820 5113
rect -786 5085 -758 5113
rect -724 5085 -696 5113
rect -910 5023 -882 5051
rect -848 5023 -820 5051
rect -786 5023 -758 5051
rect -724 5023 -696 5051
rect -910 4961 -882 4989
rect -848 4961 -820 4989
rect -786 4961 -758 4989
rect -724 4961 -696 4989
rect -430 298578 -402 298606
rect -368 298578 -340 298606
rect -306 298578 -278 298606
rect -244 298578 -216 298606
rect -430 298516 -402 298544
rect -368 298516 -340 298544
rect -306 298516 -278 298544
rect -244 298516 -216 298544
rect -430 298454 -402 298482
rect -368 298454 -340 298482
rect -306 298454 -278 298482
rect -244 298454 -216 298482
rect -430 298392 -402 298420
rect -368 298392 -340 298420
rect -306 298392 -278 298420
rect -244 298392 -216 298420
rect -430 290147 -402 290175
rect -368 290147 -340 290175
rect -306 290147 -278 290175
rect -244 290147 -216 290175
rect -430 290085 -402 290113
rect -368 290085 -340 290113
rect -306 290085 -278 290113
rect -244 290085 -216 290113
rect -430 290023 -402 290051
rect -368 290023 -340 290051
rect -306 290023 -278 290051
rect -244 290023 -216 290051
rect -430 289961 -402 289989
rect -368 289961 -340 289989
rect -306 289961 -278 289989
rect -244 289961 -216 289989
rect 2757 298578 2785 298606
rect 2819 298578 2847 298606
rect 2881 298578 2909 298606
rect 2943 298578 2971 298606
rect 2757 298516 2785 298544
rect 2819 298516 2847 298544
rect 2881 298516 2909 298544
rect 2943 298516 2971 298544
rect 2757 298454 2785 298482
rect 2819 298454 2847 298482
rect 2881 298454 2909 298482
rect 2943 298454 2971 298482
rect 2757 298392 2785 298420
rect 2819 298392 2847 298420
rect 2881 298392 2909 298420
rect 2943 298392 2971 298420
rect 4617 299058 4645 299086
rect 4679 299058 4707 299086
rect 4741 299058 4769 299086
rect 4803 299058 4831 299086
rect 4617 298996 4645 299024
rect 4679 298996 4707 299024
rect 4741 298996 4769 299024
rect 4803 298996 4831 299024
rect 4617 298934 4645 298962
rect 4679 298934 4707 298962
rect 4741 298934 4769 298962
rect 4803 298934 4831 298962
rect 4617 298872 4645 298900
rect 4679 298872 4707 298900
rect 4741 298872 4769 298900
rect 4803 298872 4831 298900
rect 2757 290147 2785 290175
rect 2819 290147 2847 290175
rect 2881 290147 2909 290175
rect 2943 290147 2971 290175
rect 2757 290085 2785 290113
rect 2819 290085 2847 290113
rect 2881 290085 2909 290113
rect 2943 290085 2971 290113
rect 2757 290023 2785 290051
rect 2819 290023 2847 290051
rect 2881 290023 2909 290051
rect 2943 290023 2971 290051
rect 2757 289961 2785 289989
rect 2819 289961 2847 289989
rect 2881 289961 2909 289989
rect 2943 289961 2971 289989
rect -430 281147 -402 281175
rect -368 281147 -340 281175
rect -306 281147 -278 281175
rect -244 281147 -216 281175
rect -430 281085 -402 281113
rect -368 281085 -340 281113
rect -306 281085 -278 281113
rect -244 281085 -216 281113
rect -430 281023 -402 281051
rect -368 281023 -340 281051
rect -306 281023 -278 281051
rect -244 281023 -216 281051
rect -430 280961 -402 280989
rect -368 280961 -340 280989
rect -306 280961 -278 280989
rect -244 280961 -216 280989
rect -430 272147 -402 272175
rect -368 272147 -340 272175
rect -306 272147 -278 272175
rect -244 272147 -216 272175
rect -430 272085 -402 272113
rect -368 272085 -340 272113
rect -306 272085 -278 272113
rect -244 272085 -216 272113
rect -430 272023 -402 272051
rect -368 272023 -340 272051
rect -306 272023 -278 272051
rect -244 272023 -216 272051
rect -430 271961 -402 271989
rect -368 271961 -340 271989
rect -306 271961 -278 271989
rect -244 271961 -216 271989
rect -430 263147 -402 263175
rect -368 263147 -340 263175
rect -306 263147 -278 263175
rect -244 263147 -216 263175
rect -430 263085 -402 263113
rect -368 263085 -340 263113
rect -306 263085 -278 263113
rect -244 263085 -216 263113
rect -430 263023 -402 263051
rect -368 263023 -340 263051
rect -306 263023 -278 263051
rect -244 263023 -216 263051
rect -430 262961 -402 262989
rect -368 262961 -340 262989
rect -306 262961 -278 262989
rect -244 262961 -216 262989
rect -430 254147 -402 254175
rect -368 254147 -340 254175
rect -306 254147 -278 254175
rect -244 254147 -216 254175
rect -430 254085 -402 254113
rect -368 254085 -340 254113
rect -306 254085 -278 254113
rect -244 254085 -216 254113
rect -430 254023 -402 254051
rect -368 254023 -340 254051
rect -306 254023 -278 254051
rect -244 254023 -216 254051
rect -430 253961 -402 253989
rect -368 253961 -340 253989
rect -306 253961 -278 253989
rect -244 253961 -216 253989
rect -430 245147 -402 245175
rect -368 245147 -340 245175
rect -306 245147 -278 245175
rect -244 245147 -216 245175
rect -430 245085 -402 245113
rect -368 245085 -340 245113
rect -306 245085 -278 245113
rect -244 245085 -216 245113
rect -430 245023 -402 245051
rect -368 245023 -340 245051
rect -306 245023 -278 245051
rect -244 245023 -216 245051
rect -430 244961 -402 244989
rect -368 244961 -340 244989
rect -306 244961 -278 244989
rect -244 244961 -216 244989
rect -430 236147 -402 236175
rect -368 236147 -340 236175
rect -306 236147 -278 236175
rect -244 236147 -216 236175
rect -430 236085 -402 236113
rect -368 236085 -340 236113
rect -306 236085 -278 236113
rect -244 236085 -216 236113
rect -430 236023 -402 236051
rect -368 236023 -340 236051
rect -306 236023 -278 236051
rect -244 236023 -216 236051
rect -430 235961 -402 235989
rect -368 235961 -340 235989
rect -306 235961 -278 235989
rect -244 235961 -216 235989
rect -430 227147 -402 227175
rect -368 227147 -340 227175
rect -306 227147 -278 227175
rect -244 227147 -216 227175
rect -430 227085 -402 227113
rect -368 227085 -340 227113
rect -306 227085 -278 227113
rect -244 227085 -216 227113
rect -430 227023 -402 227051
rect -368 227023 -340 227051
rect -306 227023 -278 227051
rect -244 227023 -216 227051
rect -430 226961 -402 226989
rect -368 226961 -340 226989
rect -306 226961 -278 226989
rect -244 226961 -216 226989
rect -430 218147 -402 218175
rect -368 218147 -340 218175
rect -306 218147 -278 218175
rect -244 218147 -216 218175
rect -430 218085 -402 218113
rect -368 218085 -340 218113
rect -306 218085 -278 218113
rect -244 218085 -216 218113
rect -430 218023 -402 218051
rect -368 218023 -340 218051
rect -306 218023 -278 218051
rect -244 218023 -216 218051
rect -430 217961 -402 217989
rect -368 217961 -340 217989
rect -306 217961 -278 217989
rect -244 217961 -216 217989
rect -430 209147 -402 209175
rect -368 209147 -340 209175
rect -306 209147 -278 209175
rect -244 209147 -216 209175
rect -430 209085 -402 209113
rect -368 209085 -340 209113
rect -306 209085 -278 209113
rect -244 209085 -216 209113
rect -430 209023 -402 209051
rect -368 209023 -340 209051
rect -306 209023 -278 209051
rect -244 209023 -216 209051
rect -430 208961 -402 208989
rect -368 208961 -340 208989
rect -306 208961 -278 208989
rect -244 208961 -216 208989
rect -430 200147 -402 200175
rect -368 200147 -340 200175
rect -306 200147 -278 200175
rect -244 200147 -216 200175
rect -430 200085 -402 200113
rect -368 200085 -340 200113
rect -306 200085 -278 200113
rect -244 200085 -216 200113
rect -430 200023 -402 200051
rect -368 200023 -340 200051
rect -306 200023 -278 200051
rect -244 200023 -216 200051
rect -430 199961 -402 199989
rect -368 199961 -340 199989
rect -306 199961 -278 199989
rect -244 199961 -216 199989
rect -430 191147 -402 191175
rect -368 191147 -340 191175
rect -306 191147 -278 191175
rect -244 191147 -216 191175
rect -430 191085 -402 191113
rect -368 191085 -340 191113
rect -306 191085 -278 191113
rect -244 191085 -216 191113
rect -430 191023 -402 191051
rect -368 191023 -340 191051
rect -306 191023 -278 191051
rect -244 191023 -216 191051
rect -430 190961 -402 190989
rect -368 190961 -340 190989
rect -306 190961 -278 190989
rect -244 190961 -216 190989
rect -430 182147 -402 182175
rect -368 182147 -340 182175
rect -306 182147 -278 182175
rect -244 182147 -216 182175
rect -430 182085 -402 182113
rect -368 182085 -340 182113
rect -306 182085 -278 182113
rect -244 182085 -216 182113
rect -430 182023 -402 182051
rect -368 182023 -340 182051
rect -306 182023 -278 182051
rect -244 182023 -216 182051
rect -430 181961 -402 181989
rect -368 181961 -340 181989
rect -306 181961 -278 181989
rect -244 181961 -216 181989
rect -430 173147 -402 173175
rect -368 173147 -340 173175
rect -306 173147 -278 173175
rect -244 173147 -216 173175
rect -430 173085 -402 173113
rect -368 173085 -340 173113
rect -306 173085 -278 173113
rect -244 173085 -216 173113
rect -430 173023 -402 173051
rect -368 173023 -340 173051
rect -306 173023 -278 173051
rect -244 173023 -216 173051
rect -430 172961 -402 172989
rect -368 172961 -340 172989
rect -306 172961 -278 172989
rect -244 172961 -216 172989
rect -430 164147 -402 164175
rect -368 164147 -340 164175
rect -306 164147 -278 164175
rect -244 164147 -216 164175
rect -430 164085 -402 164113
rect -368 164085 -340 164113
rect -306 164085 -278 164113
rect -244 164085 -216 164113
rect -430 164023 -402 164051
rect -368 164023 -340 164051
rect -306 164023 -278 164051
rect -244 164023 -216 164051
rect -430 163961 -402 163989
rect -368 163961 -340 163989
rect -306 163961 -278 163989
rect -244 163961 -216 163989
rect 2757 281147 2785 281175
rect 2819 281147 2847 281175
rect 2881 281147 2909 281175
rect 2943 281147 2971 281175
rect 2757 281085 2785 281113
rect 2819 281085 2847 281113
rect 2881 281085 2909 281113
rect 2943 281085 2971 281113
rect 2757 281023 2785 281051
rect 2819 281023 2847 281051
rect 2881 281023 2909 281051
rect 2943 281023 2971 281051
rect 2757 280961 2785 280989
rect 2819 280961 2847 280989
rect 2881 280961 2909 280989
rect 2943 280961 2971 280989
rect 2757 272147 2785 272175
rect 2819 272147 2847 272175
rect 2881 272147 2909 272175
rect 2943 272147 2971 272175
rect 2757 272085 2785 272113
rect 2819 272085 2847 272113
rect 2881 272085 2909 272113
rect 2943 272085 2971 272113
rect 2757 272023 2785 272051
rect 2819 272023 2847 272051
rect 2881 272023 2909 272051
rect 2943 272023 2971 272051
rect 2757 271961 2785 271989
rect 2819 271961 2847 271989
rect 2881 271961 2909 271989
rect 2943 271961 2971 271989
rect -430 155147 -402 155175
rect -368 155147 -340 155175
rect -306 155147 -278 155175
rect -244 155147 -216 155175
rect -430 155085 -402 155113
rect -368 155085 -340 155113
rect -306 155085 -278 155113
rect -244 155085 -216 155113
rect -430 155023 -402 155051
rect -368 155023 -340 155051
rect -306 155023 -278 155051
rect -244 155023 -216 155051
rect -430 154961 -402 154989
rect -368 154961 -340 154989
rect -306 154961 -278 154989
rect -244 154961 -216 154989
rect 2757 263147 2785 263175
rect 2819 263147 2847 263175
rect 2881 263147 2909 263175
rect 2943 263147 2971 263175
rect 2757 263085 2785 263113
rect 2819 263085 2847 263113
rect 2881 263085 2909 263113
rect 2943 263085 2971 263113
rect 2757 263023 2785 263051
rect 2819 263023 2847 263051
rect 2881 263023 2909 263051
rect 2943 263023 2971 263051
rect 2757 262961 2785 262989
rect 2819 262961 2847 262989
rect 2881 262961 2909 262989
rect 2943 262961 2971 262989
rect 2757 254147 2785 254175
rect 2819 254147 2847 254175
rect 2881 254147 2909 254175
rect 2943 254147 2971 254175
rect 2757 254085 2785 254113
rect 2819 254085 2847 254113
rect 2881 254085 2909 254113
rect 2943 254085 2971 254113
rect 2757 254023 2785 254051
rect 2819 254023 2847 254051
rect 2881 254023 2909 254051
rect 2943 254023 2971 254051
rect 2757 253961 2785 253989
rect 2819 253961 2847 253989
rect 2881 253961 2909 253989
rect 2943 253961 2971 253989
rect 2757 245147 2785 245175
rect 2819 245147 2847 245175
rect 2881 245147 2909 245175
rect 2943 245147 2971 245175
rect 2757 245085 2785 245113
rect 2819 245085 2847 245113
rect 2881 245085 2909 245113
rect 2943 245085 2971 245113
rect 2757 245023 2785 245051
rect 2819 245023 2847 245051
rect 2881 245023 2909 245051
rect 2943 245023 2971 245051
rect 2757 244961 2785 244989
rect 2819 244961 2847 244989
rect 2881 244961 2909 244989
rect 2943 244961 2971 244989
rect -430 146147 -402 146175
rect -368 146147 -340 146175
rect -306 146147 -278 146175
rect -244 146147 -216 146175
rect -430 146085 -402 146113
rect -368 146085 -340 146113
rect -306 146085 -278 146113
rect -244 146085 -216 146113
rect -430 146023 -402 146051
rect -368 146023 -340 146051
rect -306 146023 -278 146051
rect -244 146023 -216 146051
rect -430 145961 -402 145989
rect -368 145961 -340 145989
rect -306 145961 -278 145989
rect -244 145961 -216 145989
rect 2757 236147 2785 236175
rect 2819 236147 2847 236175
rect 2881 236147 2909 236175
rect 2943 236147 2971 236175
rect 2757 236085 2785 236113
rect 2819 236085 2847 236113
rect 2881 236085 2909 236113
rect 2943 236085 2971 236113
rect 2757 236023 2785 236051
rect 2819 236023 2847 236051
rect 2881 236023 2909 236051
rect 2943 236023 2971 236051
rect 2757 235961 2785 235989
rect 2819 235961 2847 235989
rect 2881 235961 2909 235989
rect 2943 235961 2971 235989
rect 2757 227147 2785 227175
rect 2819 227147 2847 227175
rect 2881 227147 2909 227175
rect 2943 227147 2971 227175
rect 2757 227085 2785 227113
rect 2819 227085 2847 227113
rect 2881 227085 2909 227113
rect 2943 227085 2971 227113
rect 2757 227023 2785 227051
rect 2819 227023 2847 227051
rect 2881 227023 2909 227051
rect 2943 227023 2971 227051
rect 2757 226961 2785 226989
rect 2819 226961 2847 226989
rect 2881 226961 2909 226989
rect 2943 226961 2971 226989
rect 2757 218147 2785 218175
rect 2819 218147 2847 218175
rect 2881 218147 2909 218175
rect 2943 218147 2971 218175
rect 2757 218085 2785 218113
rect 2819 218085 2847 218113
rect 2881 218085 2909 218113
rect 2943 218085 2971 218113
rect 2757 218023 2785 218051
rect 2819 218023 2847 218051
rect 2881 218023 2909 218051
rect 2943 218023 2971 218051
rect 2757 217961 2785 217989
rect 2819 217961 2847 217989
rect 2881 217961 2909 217989
rect 2943 217961 2971 217989
rect 2757 209147 2785 209175
rect 2819 209147 2847 209175
rect 2881 209147 2909 209175
rect 2943 209147 2971 209175
rect 2757 209085 2785 209113
rect 2819 209085 2847 209113
rect 2881 209085 2909 209113
rect 2943 209085 2971 209113
rect 2757 209023 2785 209051
rect 2819 209023 2847 209051
rect 2881 209023 2909 209051
rect 2943 209023 2971 209051
rect 2757 208961 2785 208989
rect 2819 208961 2847 208989
rect 2881 208961 2909 208989
rect 2943 208961 2971 208989
rect 2757 200147 2785 200175
rect 2819 200147 2847 200175
rect 2881 200147 2909 200175
rect 2943 200147 2971 200175
rect 2757 200085 2785 200113
rect 2819 200085 2847 200113
rect 2881 200085 2909 200113
rect 2943 200085 2971 200113
rect 2757 200023 2785 200051
rect 2819 200023 2847 200051
rect 2881 200023 2909 200051
rect 2943 200023 2971 200051
rect 2757 199961 2785 199989
rect 2819 199961 2847 199989
rect 2881 199961 2909 199989
rect 2943 199961 2971 199989
rect 2757 191147 2785 191175
rect 2819 191147 2847 191175
rect 2881 191147 2909 191175
rect 2943 191147 2971 191175
rect 2757 191085 2785 191113
rect 2819 191085 2847 191113
rect 2881 191085 2909 191113
rect 2943 191085 2971 191113
rect 2757 191023 2785 191051
rect 2819 191023 2847 191051
rect 2881 191023 2909 191051
rect 2943 191023 2971 191051
rect 2757 190961 2785 190989
rect 2819 190961 2847 190989
rect 2881 190961 2909 190989
rect 2943 190961 2971 190989
rect 2757 182147 2785 182175
rect 2819 182147 2847 182175
rect 2881 182147 2909 182175
rect 2943 182147 2971 182175
rect 2757 182085 2785 182113
rect 2819 182085 2847 182113
rect 2881 182085 2909 182113
rect 2943 182085 2971 182113
rect 2757 182023 2785 182051
rect 2819 182023 2847 182051
rect 2881 182023 2909 182051
rect 2943 182023 2971 182051
rect 2757 181961 2785 181989
rect 2819 181961 2847 181989
rect 2881 181961 2909 181989
rect 2943 181961 2971 181989
rect 2757 173147 2785 173175
rect 2819 173147 2847 173175
rect 2881 173147 2909 173175
rect 2943 173147 2971 173175
rect 2757 173085 2785 173113
rect 2819 173085 2847 173113
rect 2881 173085 2909 173113
rect 2943 173085 2971 173113
rect 2757 173023 2785 173051
rect 2819 173023 2847 173051
rect 2881 173023 2909 173051
rect 2943 173023 2971 173051
rect 2757 172961 2785 172989
rect 2819 172961 2847 172989
rect 2881 172961 2909 172989
rect 2943 172961 2971 172989
rect 2757 164147 2785 164175
rect 2819 164147 2847 164175
rect 2881 164147 2909 164175
rect 2943 164147 2971 164175
rect 2757 164085 2785 164113
rect 2819 164085 2847 164113
rect 2881 164085 2909 164113
rect 2943 164085 2971 164113
rect 2757 164023 2785 164051
rect 2819 164023 2847 164051
rect 2881 164023 2909 164051
rect 2943 164023 2971 164051
rect 2757 163961 2785 163989
rect 2819 163961 2847 163989
rect 2881 163961 2909 163989
rect 2943 163961 2971 163989
rect 2757 155147 2785 155175
rect 2819 155147 2847 155175
rect 2881 155147 2909 155175
rect 2943 155147 2971 155175
rect 2757 155085 2785 155113
rect 2819 155085 2847 155113
rect 2881 155085 2909 155113
rect 2943 155085 2971 155113
rect 2757 155023 2785 155051
rect 2819 155023 2847 155051
rect 2881 155023 2909 155051
rect 2943 155023 2971 155051
rect 2757 154961 2785 154989
rect 2819 154961 2847 154989
rect 2881 154961 2909 154989
rect 2943 154961 2971 154989
rect 4617 293147 4645 293175
rect 4679 293147 4707 293175
rect 4741 293147 4769 293175
rect 4803 293147 4831 293175
rect 4617 293085 4645 293113
rect 4679 293085 4707 293113
rect 4741 293085 4769 293113
rect 4803 293085 4831 293113
rect 4617 293023 4645 293051
rect 4679 293023 4707 293051
rect 4741 293023 4769 293051
rect 4803 293023 4831 293051
rect 4617 292961 4645 292989
rect 4679 292961 4707 292989
rect 4741 292961 4769 292989
rect 4803 292961 4831 292989
rect 4617 284147 4645 284175
rect 4679 284147 4707 284175
rect 4741 284147 4769 284175
rect 4803 284147 4831 284175
rect 4617 284085 4645 284113
rect 4679 284085 4707 284113
rect 4741 284085 4769 284113
rect 4803 284085 4831 284113
rect 4617 284023 4645 284051
rect 4679 284023 4707 284051
rect 4741 284023 4769 284051
rect 4803 284023 4831 284051
rect 4617 283961 4645 283989
rect 4679 283961 4707 283989
rect 4741 283961 4769 283989
rect 4803 283961 4831 283989
rect 18117 298578 18145 298606
rect 18179 298578 18207 298606
rect 18241 298578 18269 298606
rect 18303 298578 18331 298606
rect 18117 298516 18145 298544
rect 18179 298516 18207 298544
rect 18241 298516 18269 298544
rect 18303 298516 18331 298544
rect 18117 298454 18145 298482
rect 18179 298454 18207 298482
rect 18241 298454 18269 298482
rect 18303 298454 18331 298482
rect 18117 298392 18145 298420
rect 18179 298392 18207 298420
rect 18241 298392 18269 298420
rect 18303 298392 18331 298420
rect 18117 290147 18145 290175
rect 18179 290147 18207 290175
rect 18241 290147 18269 290175
rect 18303 290147 18331 290175
rect 18117 290085 18145 290113
rect 18179 290085 18207 290113
rect 18241 290085 18269 290113
rect 18303 290085 18331 290113
rect 18117 290023 18145 290051
rect 18179 290023 18207 290051
rect 18241 290023 18269 290051
rect 18303 290023 18331 290051
rect 18117 289961 18145 289989
rect 18179 289961 18207 289989
rect 18241 289961 18269 289989
rect 18303 289961 18331 289989
rect 18117 281147 18145 281175
rect 18179 281147 18207 281175
rect 18241 281147 18269 281175
rect 18303 281147 18331 281175
rect 18117 281085 18145 281113
rect 18179 281085 18207 281113
rect 18241 281085 18269 281113
rect 18303 281085 18331 281113
rect 18117 281023 18145 281051
rect 18179 281023 18207 281051
rect 18241 281023 18269 281051
rect 18303 281023 18331 281051
rect 18117 280961 18145 280989
rect 18179 280961 18207 280989
rect 18241 280961 18269 280989
rect 18303 280961 18331 280989
rect 4617 275147 4645 275175
rect 4679 275147 4707 275175
rect 4741 275147 4769 275175
rect 4803 275147 4831 275175
rect 4617 275085 4645 275113
rect 4679 275085 4707 275113
rect 4741 275085 4769 275113
rect 4803 275085 4831 275113
rect 4617 275023 4645 275051
rect 4679 275023 4707 275051
rect 4741 275023 4769 275051
rect 4803 275023 4831 275051
rect 4617 274961 4645 274989
rect 4679 274961 4707 274989
rect 4741 274961 4769 274989
rect 4803 274961 4831 274989
rect 4617 266147 4645 266175
rect 4679 266147 4707 266175
rect 4741 266147 4769 266175
rect 4803 266147 4831 266175
rect 4617 266085 4645 266113
rect 4679 266085 4707 266113
rect 4741 266085 4769 266113
rect 4803 266085 4831 266113
rect 4617 266023 4645 266051
rect 4679 266023 4707 266051
rect 4741 266023 4769 266051
rect 4803 266023 4831 266051
rect 4617 265961 4645 265989
rect 4679 265961 4707 265989
rect 4741 265961 4769 265989
rect 4803 265961 4831 265989
rect 4617 257147 4645 257175
rect 4679 257147 4707 257175
rect 4741 257147 4769 257175
rect 4803 257147 4831 257175
rect 4617 257085 4645 257113
rect 4679 257085 4707 257113
rect 4741 257085 4769 257113
rect 4803 257085 4831 257113
rect 4617 257023 4645 257051
rect 4679 257023 4707 257051
rect 4741 257023 4769 257051
rect 4803 257023 4831 257051
rect 4617 256961 4645 256989
rect 4679 256961 4707 256989
rect 4741 256961 4769 256989
rect 4803 256961 4831 256989
rect 4617 248147 4645 248175
rect 4679 248147 4707 248175
rect 4741 248147 4769 248175
rect 4803 248147 4831 248175
rect 4617 248085 4645 248113
rect 4679 248085 4707 248113
rect 4741 248085 4769 248113
rect 4803 248085 4831 248113
rect 4617 248023 4645 248051
rect 4679 248023 4707 248051
rect 4741 248023 4769 248051
rect 4803 248023 4831 248051
rect 4617 247961 4645 247989
rect 4679 247961 4707 247989
rect 4741 247961 4769 247989
rect 4803 247961 4831 247989
rect 4617 239147 4645 239175
rect 4679 239147 4707 239175
rect 4741 239147 4769 239175
rect 4803 239147 4831 239175
rect 4617 239085 4645 239113
rect 4679 239085 4707 239113
rect 4741 239085 4769 239113
rect 4803 239085 4831 239113
rect 4617 239023 4645 239051
rect 4679 239023 4707 239051
rect 4741 239023 4769 239051
rect 4803 239023 4831 239051
rect 4617 238961 4645 238989
rect 4679 238961 4707 238989
rect 4741 238961 4769 238989
rect 4803 238961 4831 238989
rect 4617 230147 4645 230175
rect 4679 230147 4707 230175
rect 4741 230147 4769 230175
rect 4803 230147 4831 230175
rect 4617 230085 4645 230113
rect 4679 230085 4707 230113
rect 4741 230085 4769 230113
rect 4803 230085 4831 230113
rect 4617 230023 4645 230051
rect 4679 230023 4707 230051
rect 4741 230023 4769 230051
rect 4803 230023 4831 230051
rect 4617 229961 4645 229989
rect 4679 229961 4707 229989
rect 4741 229961 4769 229989
rect 4803 229961 4831 229989
rect 4617 221147 4645 221175
rect 4679 221147 4707 221175
rect 4741 221147 4769 221175
rect 4803 221147 4831 221175
rect 4617 221085 4645 221113
rect 4679 221085 4707 221113
rect 4741 221085 4769 221113
rect 4803 221085 4831 221113
rect 4617 221023 4645 221051
rect 4679 221023 4707 221051
rect 4741 221023 4769 221051
rect 4803 221023 4831 221051
rect 4617 220961 4645 220989
rect 4679 220961 4707 220989
rect 4741 220961 4769 220989
rect 4803 220961 4831 220989
rect 4617 212147 4645 212175
rect 4679 212147 4707 212175
rect 4741 212147 4769 212175
rect 4803 212147 4831 212175
rect 4617 212085 4645 212113
rect 4679 212085 4707 212113
rect 4741 212085 4769 212113
rect 4803 212085 4831 212113
rect 4617 212023 4645 212051
rect 4679 212023 4707 212051
rect 4741 212023 4769 212051
rect 4803 212023 4831 212051
rect 4617 211961 4645 211989
rect 4679 211961 4707 211989
rect 4741 211961 4769 211989
rect 4803 211961 4831 211989
rect 4617 203147 4645 203175
rect 4679 203147 4707 203175
rect 4741 203147 4769 203175
rect 4803 203147 4831 203175
rect 4617 203085 4645 203113
rect 4679 203085 4707 203113
rect 4741 203085 4769 203113
rect 4803 203085 4831 203113
rect 4617 203023 4645 203051
rect 4679 203023 4707 203051
rect 4741 203023 4769 203051
rect 4803 203023 4831 203051
rect 4617 202961 4645 202989
rect 4679 202961 4707 202989
rect 4741 202961 4769 202989
rect 4803 202961 4831 202989
rect 4617 194147 4645 194175
rect 4679 194147 4707 194175
rect 4741 194147 4769 194175
rect 4803 194147 4831 194175
rect 4617 194085 4645 194113
rect 4679 194085 4707 194113
rect 4741 194085 4769 194113
rect 4803 194085 4831 194113
rect 4617 194023 4645 194051
rect 4679 194023 4707 194051
rect 4741 194023 4769 194051
rect 4803 194023 4831 194051
rect 4617 193961 4645 193989
rect 4679 193961 4707 193989
rect 4741 193961 4769 193989
rect 4803 193961 4831 193989
rect 4617 185147 4645 185175
rect 4679 185147 4707 185175
rect 4741 185147 4769 185175
rect 4803 185147 4831 185175
rect 4617 185085 4645 185113
rect 4679 185085 4707 185113
rect 4741 185085 4769 185113
rect 4803 185085 4831 185113
rect 4617 185023 4645 185051
rect 4679 185023 4707 185051
rect 4741 185023 4769 185051
rect 4803 185023 4831 185051
rect 4617 184961 4645 184989
rect 4679 184961 4707 184989
rect 4741 184961 4769 184989
rect 4803 184961 4831 184989
rect 4617 176147 4645 176175
rect 4679 176147 4707 176175
rect 4741 176147 4769 176175
rect 4803 176147 4831 176175
rect 4617 176085 4645 176113
rect 4679 176085 4707 176113
rect 4741 176085 4769 176113
rect 4803 176085 4831 176113
rect 4617 176023 4645 176051
rect 4679 176023 4707 176051
rect 4741 176023 4769 176051
rect 4803 176023 4831 176051
rect 4617 175961 4645 175989
rect 4679 175961 4707 175989
rect 4741 175961 4769 175989
rect 4803 175961 4831 175989
rect 4617 167147 4645 167175
rect 4679 167147 4707 167175
rect 4741 167147 4769 167175
rect 4803 167147 4831 167175
rect 4617 167085 4645 167113
rect 4679 167085 4707 167113
rect 4741 167085 4769 167113
rect 4803 167085 4831 167113
rect 4617 167023 4645 167051
rect 4679 167023 4707 167051
rect 4741 167023 4769 167051
rect 4803 167023 4831 167051
rect 4617 166961 4645 166989
rect 4679 166961 4707 166989
rect 4741 166961 4769 166989
rect 4803 166961 4831 166989
rect 2757 146147 2785 146175
rect 2819 146147 2847 146175
rect 2881 146147 2909 146175
rect 2943 146147 2971 146175
rect 2757 146085 2785 146113
rect 2819 146085 2847 146113
rect 2881 146085 2909 146113
rect 2943 146085 2971 146113
rect 2757 146023 2785 146051
rect 2819 146023 2847 146051
rect 2881 146023 2909 146051
rect 2943 146023 2971 146051
rect 4617 158147 4645 158175
rect 4679 158147 4707 158175
rect 4741 158147 4769 158175
rect 4803 158147 4831 158175
rect 4617 158085 4645 158113
rect 4679 158085 4707 158113
rect 4741 158085 4769 158113
rect 4803 158085 4831 158113
rect 4617 158023 4645 158051
rect 4679 158023 4707 158051
rect 4741 158023 4769 158051
rect 4803 158023 4831 158051
rect 4617 157961 4645 157989
rect 4679 157961 4707 157989
rect 4741 157961 4769 157989
rect 4803 157961 4831 157989
rect 4617 149147 4645 149175
rect 4679 149147 4707 149175
rect 4741 149147 4769 149175
rect 4803 149147 4831 149175
rect 4617 149085 4645 149113
rect 4679 149085 4707 149113
rect 4741 149085 4769 149113
rect 4803 149085 4831 149113
rect 4617 149023 4645 149051
rect 4679 149023 4707 149051
rect 4741 149023 4769 149051
rect 4803 149023 4831 149051
rect 4617 148961 4645 148989
rect 4679 148961 4707 148989
rect 4741 148961 4769 148989
rect 4803 148961 4831 148989
rect 2757 145961 2785 145989
rect 2819 145961 2847 145989
rect 2881 145961 2909 145989
rect 2943 145961 2971 145989
rect -430 137147 -402 137175
rect -368 137147 -340 137175
rect -306 137147 -278 137175
rect -244 137147 -216 137175
rect -430 137085 -402 137113
rect -368 137085 -340 137113
rect -306 137085 -278 137113
rect -244 137085 -216 137113
rect -430 137023 -402 137051
rect -368 137023 -340 137051
rect -306 137023 -278 137051
rect -244 137023 -216 137051
rect -430 136961 -402 136989
rect -368 136961 -340 136989
rect -306 136961 -278 136989
rect -244 136961 -216 136989
rect -430 128147 -402 128175
rect -368 128147 -340 128175
rect -306 128147 -278 128175
rect -244 128147 -216 128175
rect -430 128085 -402 128113
rect -368 128085 -340 128113
rect -306 128085 -278 128113
rect -244 128085 -216 128113
rect -430 128023 -402 128051
rect -368 128023 -340 128051
rect -306 128023 -278 128051
rect -244 128023 -216 128051
rect -430 127961 -402 127989
rect -368 127961 -340 127989
rect -306 127961 -278 127989
rect -244 127961 -216 127989
rect -430 119147 -402 119175
rect -368 119147 -340 119175
rect -306 119147 -278 119175
rect -244 119147 -216 119175
rect -430 119085 -402 119113
rect -368 119085 -340 119113
rect -306 119085 -278 119113
rect -244 119085 -216 119113
rect -430 119023 -402 119051
rect -368 119023 -340 119051
rect -306 119023 -278 119051
rect -244 119023 -216 119051
rect -430 118961 -402 118989
rect -368 118961 -340 118989
rect -306 118961 -278 118989
rect -244 118961 -216 118989
rect -430 110147 -402 110175
rect -368 110147 -340 110175
rect -306 110147 -278 110175
rect -244 110147 -216 110175
rect -430 110085 -402 110113
rect -368 110085 -340 110113
rect -306 110085 -278 110113
rect -244 110085 -216 110113
rect -430 110023 -402 110051
rect -368 110023 -340 110051
rect -306 110023 -278 110051
rect -244 110023 -216 110051
rect -430 109961 -402 109989
rect -368 109961 -340 109989
rect -306 109961 -278 109989
rect -244 109961 -216 109989
rect -430 101147 -402 101175
rect -368 101147 -340 101175
rect -306 101147 -278 101175
rect -244 101147 -216 101175
rect -430 101085 -402 101113
rect -368 101085 -340 101113
rect -306 101085 -278 101113
rect -244 101085 -216 101113
rect -430 101023 -402 101051
rect -368 101023 -340 101051
rect -306 101023 -278 101051
rect -244 101023 -216 101051
rect -430 100961 -402 100989
rect -368 100961 -340 100989
rect -306 100961 -278 100989
rect -244 100961 -216 100989
rect -430 92147 -402 92175
rect -368 92147 -340 92175
rect -306 92147 -278 92175
rect -244 92147 -216 92175
rect -430 92085 -402 92113
rect -368 92085 -340 92113
rect -306 92085 -278 92113
rect -244 92085 -216 92113
rect -430 92023 -402 92051
rect -368 92023 -340 92051
rect -306 92023 -278 92051
rect -244 92023 -216 92051
rect -430 91961 -402 91989
rect -368 91961 -340 91989
rect -306 91961 -278 91989
rect -244 91961 -216 91989
rect -430 83147 -402 83175
rect -368 83147 -340 83175
rect -306 83147 -278 83175
rect -244 83147 -216 83175
rect -430 83085 -402 83113
rect -368 83085 -340 83113
rect -306 83085 -278 83113
rect -244 83085 -216 83113
rect -430 83023 -402 83051
rect -368 83023 -340 83051
rect -306 83023 -278 83051
rect -244 83023 -216 83051
rect -430 82961 -402 82989
rect -368 82961 -340 82989
rect -306 82961 -278 82989
rect -244 82961 -216 82989
rect -430 74147 -402 74175
rect -368 74147 -340 74175
rect -306 74147 -278 74175
rect -244 74147 -216 74175
rect -430 74085 -402 74113
rect -368 74085 -340 74113
rect -306 74085 -278 74113
rect -244 74085 -216 74113
rect -430 74023 -402 74051
rect -368 74023 -340 74051
rect -306 74023 -278 74051
rect -244 74023 -216 74051
rect -430 73961 -402 73989
rect -368 73961 -340 73989
rect -306 73961 -278 73989
rect -244 73961 -216 73989
rect -430 65147 -402 65175
rect -368 65147 -340 65175
rect -306 65147 -278 65175
rect -244 65147 -216 65175
rect -430 65085 -402 65113
rect -368 65085 -340 65113
rect -306 65085 -278 65113
rect -244 65085 -216 65113
rect -430 65023 -402 65051
rect -368 65023 -340 65051
rect -306 65023 -278 65051
rect -244 65023 -216 65051
rect -430 64961 -402 64989
rect -368 64961 -340 64989
rect -306 64961 -278 64989
rect -244 64961 -216 64989
rect -430 56147 -402 56175
rect -368 56147 -340 56175
rect -306 56147 -278 56175
rect -244 56147 -216 56175
rect -430 56085 -402 56113
rect -368 56085 -340 56113
rect -306 56085 -278 56113
rect -244 56085 -216 56113
rect -430 56023 -402 56051
rect -368 56023 -340 56051
rect -306 56023 -278 56051
rect -244 56023 -216 56051
rect -430 55961 -402 55989
rect -368 55961 -340 55989
rect -306 55961 -278 55989
rect -244 55961 -216 55989
rect -430 47147 -402 47175
rect -368 47147 -340 47175
rect -306 47147 -278 47175
rect -244 47147 -216 47175
rect -430 47085 -402 47113
rect -368 47085 -340 47113
rect -306 47085 -278 47113
rect -244 47085 -216 47113
rect -430 47023 -402 47051
rect -368 47023 -340 47051
rect -306 47023 -278 47051
rect -244 47023 -216 47051
rect -430 46961 -402 46989
rect -368 46961 -340 46989
rect -306 46961 -278 46989
rect -244 46961 -216 46989
rect -430 38147 -402 38175
rect -368 38147 -340 38175
rect -306 38147 -278 38175
rect -244 38147 -216 38175
rect -430 38085 -402 38113
rect -368 38085 -340 38113
rect -306 38085 -278 38113
rect -244 38085 -216 38113
rect -430 38023 -402 38051
rect -368 38023 -340 38051
rect -306 38023 -278 38051
rect -244 38023 -216 38051
rect -430 37961 -402 37989
rect -368 37961 -340 37989
rect -306 37961 -278 37989
rect -244 37961 -216 37989
rect -430 29147 -402 29175
rect -368 29147 -340 29175
rect -306 29147 -278 29175
rect -244 29147 -216 29175
rect -430 29085 -402 29113
rect -368 29085 -340 29113
rect -306 29085 -278 29113
rect -244 29085 -216 29113
rect -430 29023 -402 29051
rect -368 29023 -340 29051
rect -306 29023 -278 29051
rect -244 29023 -216 29051
rect -430 28961 -402 28989
rect -368 28961 -340 28989
rect -306 28961 -278 28989
rect -244 28961 -216 28989
rect -430 20147 -402 20175
rect -368 20147 -340 20175
rect -306 20147 -278 20175
rect -244 20147 -216 20175
rect -430 20085 -402 20113
rect -368 20085 -340 20113
rect -306 20085 -278 20113
rect -244 20085 -216 20113
rect -430 20023 -402 20051
rect -368 20023 -340 20051
rect -306 20023 -278 20051
rect -244 20023 -216 20051
rect -430 19961 -402 19989
rect -368 19961 -340 19989
rect -306 19961 -278 19989
rect -244 19961 -216 19989
rect -430 11147 -402 11175
rect -368 11147 -340 11175
rect -306 11147 -278 11175
rect -244 11147 -216 11175
rect -430 11085 -402 11113
rect -368 11085 -340 11113
rect -306 11085 -278 11113
rect -244 11085 -216 11113
rect -430 11023 -402 11051
rect -368 11023 -340 11051
rect -306 11023 -278 11051
rect -244 11023 -216 11051
rect -430 10961 -402 10989
rect -368 10961 -340 10989
rect -306 10961 -278 10989
rect -244 10961 -216 10989
rect 2757 137147 2785 137175
rect 2819 137147 2847 137175
rect 2881 137147 2909 137175
rect 2943 137147 2971 137175
rect 2757 137085 2785 137113
rect 2819 137085 2847 137113
rect 2881 137085 2909 137113
rect 2943 137085 2971 137113
rect 2757 137023 2785 137051
rect 2819 137023 2847 137051
rect 2881 137023 2909 137051
rect 2943 137023 2971 137051
rect 2757 136961 2785 136989
rect 2819 136961 2847 136989
rect 2881 136961 2909 136989
rect 2943 136961 2971 136989
rect 2757 128147 2785 128175
rect 2819 128147 2847 128175
rect 2881 128147 2909 128175
rect 2943 128147 2971 128175
rect 2757 128085 2785 128113
rect 2819 128085 2847 128113
rect 2881 128085 2909 128113
rect 2943 128085 2971 128113
rect 2757 128023 2785 128051
rect 2819 128023 2847 128051
rect 2881 128023 2909 128051
rect 2943 128023 2971 128051
rect 2757 127961 2785 127989
rect 2819 127961 2847 127989
rect 2881 127961 2909 127989
rect 2943 127961 2971 127989
rect 2757 119147 2785 119175
rect 2819 119147 2847 119175
rect 2881 119147 2909 119175
rect 2943 119147 2971 119175
rect 2757 119085 2785 119113
rect 2819 119085 2847 119113
rect 2881 119085 2909 119113
rect 2943 119085 2971 119113
rect 2757 119023 2785 119051
rect 2819 119023 2847 119051
rect 2881 119023 2909 119051
rect 2943 119023 2971 119051
rect 2757 118961 2785 118989
rect 2819 118961 2847 118989
rect 2881 118961 2909 118989
rect 2943 118961 2971 118989
rect 2757 110147 2785 110175
rect 2819 110147 2847 110175
rect 2881 110147 2909 110175
rect 2943 110147 2971 110175
rect 2757 110085 2785 110113
rect 2819 110085 2847 110113
rect 2881 110085 2909 110113
rect 2943 110085 2971 110113
rect 2757 110023 2785 110051
rect 2819 110023 2847 110051
rect 2881 110023 2909 110051
rect 2943 110023 2971 110051
rect 2757 109961 2785 109989
rect 2819 109961 2847 109989
rect 2881 109961 2909 109989
rect 2943 109961 2971 109989
rect 2757 101147 2785 101175
rect 2819 101147 2847 101175
rect 2881 101147 2909 101175
rect 2943 101147 2971 101175
rect 2757 101085 2785 101113
rect 2819 101085 2847 101113
rect 2881 101085 2909 101113
rect 2943 101085 2971 101113
rect 2757 101023 2785 101051
rect 2819 101023 2847 101051
rect 2881 101023 2909 101051
rect 2943 101023 2971 101051
rect 2757 100961 2785 100989
rect 2819 100961 2847 100989
rect 2881 100961 2909 100989
rect 2943 100961 2971 100989
rect 2757 92147 2785 92175
rect 2819 92147 2847 92175
rect 2881 92147 2909 92175
rect 2943 92147 2971 92175
rect 2757 92085 2785 92113
rect 2819 92085 2847 92113
rect 2881 92085 2909 92113
rect 2943 92085 2971 92113
rect 2757 92023 2785 92051
rect 2819 92023 2847 92051
rect 2881 92023 2909 92051
rect 2943 92023 2971 92051
rect 2757 91961 2785 91989
rect 2819 91961 2847 91989
rect 2881 91961 2909 91989
rect 2943 91961 2971 91989
rect 2757 83147 2785 83175
rect 2819 83147 2847 83175
rect 2881 83147 2909 83175
rect 2943 83147 2971 83175
rect 2757 83085 2785 83113
rect 2819 83085 2847 83113
rect 2881 83085 2909 83113
rect 2943 83085 2971 83113
rect 2757 83023 2785 83051
rect 2819 83023 2847 83051
rect 2881 83023 2909 83051
rect 2943 83023 2971 83051
rect 2757 82961 2785 82989
rect 2819 82961 2847 82989
rect 2881 82961 2909 82989
rect 2943 82961 2971 82989
rect 2757 74147 2785 74175
rect 2819 74147 2847 74175
rect 2881 74147 2909 74175
rect 2943 74147 2971 74175
rect 2757 74085 2785 74113
rect 2819 74085 2847 74113
rect 2881 74085 2909 74113
rect 2943 74085 2971 74113
rect 2757 74023 2785 74051
rect 2819 74023 2847 74051
rect 2881 74023 2909 74051
rect 2943 74023 2971 74051
rect 2757 73961 2785 73989
rect 2819 73961 2847 73989
rect 2881 73961 2909 73989
rect 2943 73961 2971 73989
rect 2757 65147 2785 65175
rect 2819 65147 2847 65175
rect 2881 65147 2909 65175
rect 2943 65147 2971 65175
rect 2757 65085 2785 65113
rect 2819 65085 2847 65113
rect 2881 65085 2909 65113
rect 2943 65085 2971 65113
rect 2757 65023 2785 65051
rect 2819 65023 2847 65051
rect 2881 65023 2909 65051
rect 2943 65023 2971 65051
rect 2757 64961 2785 64989
rect 2819 64961 2847 64989
rect 2881 64961 2909 64989
rect 2943 64961 2971 64989
rect 2757 56147 2785 56175
rect 2819 56147 2847 56175
rect 2881 56147 2909 56175
rect 2943 56147 2971 56175
rect 2757 56085 2785 56113
rect 2819 56085 2847 56113
rect 2881 56085 2909 56113
rect 2943 56085 2971 56113
rect 2757 56023 2785 56051
rect 2819 56023 2847 56051
rect 2881 56023 2909 56051
rect 2943 56023 2971 56051
rect 2757 55961 2785 55989
rect 2819 55961 2847 55989
rect 2881 55961 2909 55989
rect 2943 55961 2971 55989
rect 2757 47147 2785 47175
rect 2819 47147 2847 47175
rect 2881 47147 2909 47175
rect 2943 47147 2971 47175
rect 2757 47085 2785 47113
rect 2819 47085 2847 47113
rect 2881 47085 2909 47113
rect 2943 47085 2971 47113
rect 2757 47023 2785 47051
rect 2819 47023 2847 47051
rect 2881 47023 2909 47051
rect 2943 47023 2971 47051
rect 2757 46961 2785 46989
rect 2819 46961 2847 46989
rect 2881 46961 2909 46989
rect 2943 46961 2971 46989
rect 18117 272147 18145 272175
rect 18179 272147 18207 272175
rect 18241 272147 18269 272175
rect 18303 272147 18331 272175
rect 18117 272085 18145 272113
rect 18179 272085 18207 272113
rect 18241 272085 18269 272113
rect 18303 272085 18331 272113
rect 18117 272023 18145 272051
rect 18179 272023 18207 272051
rect 18241 272023 18269 272051
rect 18303 272023 18331 272051
rect 18117 271961 18145 271989
rect 18179 271961 18207 271989
rect 18241 271961 18269 271989
rect 18303 271961 18331 271989
rect 19977 299058 20005 299086
rect 20039 299058 20067 299086
rect 20101 299058 20129 299086
rect 20163 299058 20191 299086
rect 19977 298996 20005 299024
rect 20039 298996 20067 299024
rect 20101 298996 20129 299024
rect 20163 298996 20191 299024
rect 19977 298934 20005 298962
rect 20039 298934 20067 298962
rect 20101 298934 20129 298962
rect 20163 298934 20191 298962
rect 19977 298872 20005 298900
rect 20039 298872 20067 298900
rect 20101 298872 20129 298900
rect 20163 298872 20191 298900
rect 19977 293147 20005 293175
rect 20039 293147 20067 293175
rect 20101 293147 20129 293175
rect 20163 293147 20191 293175
rect 19977 293085 20005 293113
rect 20039 293085 20067 293113
rect 20101 293085 20129 293113
rect 20163 293085 20191 293113
rect 19977 293023 20005 293051
rect 20039 293023 20067 293051
rect 20101 293023 20129 293051
rect 20163 293023 20191 293051
rect 19977 292961 20005 292989
rect 20039 292961 20067 292989
rect 20101 292961 20129 292989
rect 20163 292961 20191 292989
rect 19977 284147 20005 284175
rect 20039 284147 20067 284175
rect 20101 284147 20129 284175
rect 20163 284147 20191 284175
rect 19977 284085 20005 284113
rect 20039 284085 20067 284113
rect 20101 284085 20129 284113
rect 20163 284085 20191 284113
rect 19977 284023 20005 284051
rect 20039 284023 20067 284051
rect 20101 284023 20129 284051
rect 20163 284023 20191 284051
rect 19977 283961 20005 283989
rect 20039 283961 20067 283989
rect 20101 283961 20129 283989
rect 20163 283961 20191 283989
rect 19977 275147 20005 275175
rect 20039 275147 20067 275175
rect 20101 275147 20129 275175
rect 20163 275147 20191 275175
rect 19977 275085 20005 275113
rect 20039 275085 20067 275113
rect 20101 275085 20129 275113
rect 20163 275085 20191 275113
rect 19977 275023 20005 275051
rect 20039 275023 20067 275051
rect 20101 275023 20129 275051
rect 20163 275023 20191 275051
rect 19977 274961 20005 274989
rect 20039 274961 20067 274989
rect 20101 274961 20129 274989
rect 20163 274961 20191 274989
rect 33477 298578 33505 298606
rect 33539 298578 33567 298606
rect 33601 298578 33629 298606
rect 33663 298578 33691 298606
rect 33477 298516 33505 298544
rect 33539 298516 33567 298544
rect 33601 298516 33629 298544
rect 33663 298516 33691 298544
rect 33477 298454 33505 298482
rect 33539 298454 33567 298482
rect 33601 298454 33629 298482
rect 33663 298454 33691 298482
rect 33477 298392 33505 298420
rect 33539 298392 33567 298420
rect 33601 298392 33629 298420
rect 33663 298392 33691 298420
rect 33477 290147 33505 290175
rect 33539 290147 33567 290175
rect 33601 290147 33629 290175
rect 33663 290147 33691 290175
rect 33477 290085 33505 290113
rect 33539 290085 33567 290113
rect 33601 290085 33629 290113
rect 33663 290085 33691 290113
rect 33477 290023 33505 290051
rect 33539 290023 33567 290051
rect 33601 290023 33629 290051
rect 33663 290023 33691 290051
rect 33477 289961 33505 289989
rect 33539 289961 33567 289989
rect 33601 289961 33629 289989
rect 33663 289961 33691 289989
rect 33477 281147 33505 281175
rect 33539 281147 33567 281175
rect 33601 281147 33629 281175
rect 33663 281147 33691 281175
rect 33477 281085 33505 281113
rect 33539 281085 33567 281113
rect 33601 281085 33629 281113
rect 33663 281085 33691 281113
rect 33477 281023 33505 281051
rect 33539 281023 33567 281051
rect 33601 281023 33629 281051
rect 33663 281023 33691 281051
rect 33477 280961 33505 280989
rect 33539 280961 33567 280989
rect 33601 280961 33629 280989
rect 33663 280961 33691 280989
rect 33477 272147 33505 272175
rect 33539 272147 33567 272175
rect 33601 272147 33629 272175
rect 33663 272147 33691 272175
rect 33477 272085 33505 272113
rect 33539 272085 33567 272113
rect 33601 272085 33629 272113
rect 33663 272085 33691 272113
rect 33477 272023 33505 272051
rect 33539 272023 33567 272051
rect 33601 272023 33629 272051
rect 33663 272023 33691 272051
rect 33477 271961 33505 271989
rect 33539 271961 33567 271989
rect 33601 271961 33629 271989
rect 33663 271961 33691 271989
rect 35337 299058 35365 299086
rect 35399 299058 35427 299086
rect 35461 299058 35489 299086
rect 35523 299058 35551 299086
rect 35337 298996 35365 299024
rect 35399 298996 35427 299024
rect 35461 298996 35489 299024
rect 35523 298996 35551 299024
rect 35337 298934 35365 298962
rect 35399 298934 35427 298962
rect 35461 298934 35489 298962
rect 35523 298934 35551 298962
rect 35337 298872 35365 298900
rect 35399 298872 35427 298900
rect 35461 298872 35489 298900
rect 35523 298872 35551 298900
rect 35337 293147 35365 293175
rect 35399 293147 35427 293175
rect 35461 293147 35489 293175
rect 35523 293147 35551 293175
rect 35337 293085 35365 293113
rect 35399 293085 35427 293113
rect 35461 293085 35489 293113
rect 35523 293085 35551 293113
rect 35337 293023 35365 293051
rect 35399 293023 35427 293051
rect 35461 293023 35489 293051
rect 35523 293023 35551 293051
rect 35337 292961 35365 292989
rect 35399 292961 35427 292989
rect 35461 292961 35489 292989
rect 35523 292961 35551 292989
rect 35337 284147 35365 284175
rect 35399 284147 35427 284175
rect 35461 284147 35489 284175
rect 35523 284147 35551 284175
rect 35337 284085 35365 284113
rect 35399 284085 35427 284113
rect 35461 284085 35489 284113
rect 35523 284085 35551 284113
rect 35337 284023 35365 284051
rect 35399 284023 35427 284051
rect 35461 284023 35489 284051
rect 35523 284023 35551 284051
rect 35337 283961 35365 283989
rect 35399 283961 35427 283989
rect 35461 283961 35489 283989
rect 35523 283961 35551 283989
rect 35337 275147 35365 275175
rect 35399 275147 35427 275175
rect 35461 275147 35489 275175
rect 35523 275147 35551 275175
rect 35337 275085 35365 275113
rect 35399 275085 35427 275113
rect 35461 275085 35489 275113
rect 35523 275085 35551 275113
rect 35337 275023 35365 275051
rect 35399 275023 35427 275051
rect 35461 275023 35489 275051
rect 35523 275023 35551 275051
rect 35337 274961 35365 274989
rect 35399 274961 35427 274989
rect 35461 274961 35489 274989
rect 35523 274961 35551 274989
rect 48837 298578 48865 298606
rect 48899 298578 48927 298606
rect 48961 298578 48989 298606
rect 49023 298578 49051 298606
rect 48837 298516 48865 298544
rect 48899 298516 48927 298544
rect 48961 298516 48989 298544
rect 49023 298516 49051 298544
rect 48837 298454 48865 298482
rect 48899 298454 48927 298482
rect 48961 298454 48989 298482
rect 49023 298454 49051 298482
rect 48837 298392 48865 298420
rect 48899 298392 48927 298420
rect 48961 298392 48989 298420
rect 49023 298392 49051 298420
rect 48837 290147 48865 290175
rect 48899 290147 48927 290175
rect 48961 290147 48989 290175
rect 49023 290147 49051 290175
rect 48837 290085 48865 290113
rect 48899 290085 48927 290113
rect 48961 290085 48989 290113
rect 49023 290085 49051 290113
rect 48837 290023 48865 290051
rect 48899 290023 48927 290051
rect 48961 290023 48989 290051
rect 49023 290023 49051 290051
rect 48837 289961 48865 289989
rect 48899 289961 48927 289989
rect 48961 289961 48989 289989
rect 49023 289961 49051 289989
rect 48837 281147 48865 281175
rect 48899 281147 48927 281175
rect 48961 281147 48989 281175
rect 49023 281147 49051 281175
rect 48837 281085 48865 281113
rect 48899 281085 48927 281113
rect 48961 281085 48989 281113
rect 49023 281085 49051 281113
rect 48837 281023 48865 281051
rect 48899 281023 48927 281051
rect 48961 281023 48989 281051
rect 49023 281023 49051 281051
rect 48837 280961 48865 280989
rect 48899 280961 48927 280989
rect 48961 280961 48989 280989
rect 49023 280961 49051 280989
rect 48837 272147 48865 272175
rect 48899 272147 48927 272175
rect 48961 272147 48989 272175
rect 49023 272147 49051 272175
rect 48837 272085 48865 272113
rect 48899 272085 48927 272113
rect 48961 272085 48989 272113
rect 49023 272085 49051 272113
rect 48837 272023 48865 272051
rect 48899 272023 48927 272051
rect 48961 272023 48989 272051
rect 49023 272023 49051 272051
rect 48837 271961 48865 271989
rect 48899 271961 48927 271989
rect 48961 271961 48989 271989
rect 49023 271961 49051 271989
rect 50697 299058 50725 299086
rect 50759 299058 50787 299086
rect 50821 299058 50849 299086
rect 50883 299058 50911 299086
rect 50697 298996 50725 299024
rect 50759 298996 50787 299024
rect 50821 298996 50849 299024
rect 50883 298996 50911 299024
rect 50697 298934 50725 298962
rect 50759 298934 50787 298962
rect 50821 298934 50849 298962
rect 50883 298934 50911 298962
rect 50697 298872 50725 298900
rect 50759 298872 50787 298900
rect 50821 298872 50849 298900
rect 50883 298872 50911 298900
rect 50697 293147 50725 293175
rect 50759 293147 50787 293175
rect 50821 293147 50849 293175
rect 50883 293147 50911 293175
rect 50697 293085 50725 293113
rect 50759 293085 50787 293113
rect 50821 293085 50849 293113
rect 50883 293085 50911 293113
rect 50697 293023 50725 293051
rect 50759 293023 50787 293051
rect 50821 293023 50849 293051
rect 50883 293023 50911 293051
rect 50697 292961 50725 292989
rect 50759 292961 50787 292989
rect 50821 292961 50849 292989
rect 50883 292961 50911 292989
rect 50697 284147 50725 284175
rect 50759 284147 50787 284175
rect 50821 284147 50849 284175
rect 50883 284147 50911 284175
rect 50697 284085 50725 284113
rect 50759 284085 50787 284113
rect 50821 284085 50849 284113
rect 50883 284085 50911 284113
rect 50697 284023 50725 284051
rect 50759 284023 50787 284051
rect 50821 284023 50849 284051
rect 50883 284023 50911 284051
rect 50697 283961 50725 283989
rect 50759 283961 50787 283989
rect 50821 283961 50849 283989
rect 50883 283961 50911 283989
rect 50697 275147 50725 275175
rect 50759 275147 50787 275175
rect 50821 275147 50849 275175
rect 50883 275147 50911 275175
rect 50697 275085 50725 275113
rect 50759 275085 50787 275113
rect 50821 275085 50849 275113
rect 50883 275085 50911 275113
rect 50697 275023 50725 275051
rect 50759 275023 50787 275051
rect 50821 275023 50849 275051
rect 50883 275023 50911 275051
rect 50697 274961 50725 274989
rect 50759 274961 50787 274989
rect 50821 274961 50849 274989
rect 50883 274961 50911 274989
rect 64197 298578 64225 298606
rect 64259 298578 64287 298606
rect 64321 298578 64349 298606
rect 64383 298578 64411 298606
rect 64197 298516 64225 298544
rect 64259 298516 64287 298544
rect 64321 298516 64349 298544
rect 64383 298516 64411 298544
rect 64197 298454 64225 298482
rect 64259 298454 64287 298482
rect 64321 298454 64349 298482
rect 64383 298454 64411 298482
rect 64197 298392 64225 298420
rect 64259 298392 64287 298420
rect 64321 298392 64349 298420
rect 64383 298392 64411 298420
rect 64197 290147 64225 290175
rect 64259 290147 64287 290175
rect 64321 290147 64349 290175
rect 64383 290147 64411 290175
rect 64197 290085 64225 290113
rect 64259 290085 64287 290113
rect 64321 290085 64349 290113
rect 64383 290085 64411 290113
rect 64197 290023 64225 290051
rect 64259 290023 64287 290051
rect 64321 290023 64349 290051
rect 64383 290023 64411 290051
rect 64197 289961 64225 289989
rect 64259 289961 64287 289989
rect 64321 289961 64349 289989
rect 64383 289961 64411 289989
rect 64197 281147 64225 281175
rect 64259 281147 64287 281175
rect 64321 281147 64349 281175
rect 64383 281147 64411 281175
rect 64197 281085 64225 281113
rect 64259 281085 64287 281113
rect 64321 281085 64349 281113
rect 64383 281085 64411 281113
rect 64197 281023 64225 281051
rect 64259 281023 64287 281051
rect 64321 281023 64349 281051
rect 64383 281023 64411 281051
rect 64197 280961 64225 280989
rect 64259 280961 64287 280989
rect 64321 280961 64349 280989
rect 64383 280961 64411 280989
rect 64197 272147 64225 272175
rect 64259 272147 64287 272175
rect 64321 272147 64349 272175
rect 64383 272147 64411 272175
rect 64197 272085 64225 272113
rect 64259 272085 64287 272113
rect 64321 272085 64349 272113
rect 64383 272085 64411 272113
rect 64197 272023 64225 272051
rect 64259 272023 64287 272051
rect 64321 272023 64349 272051
rect 64383 272023 64411 272051
rect 64197 271961 64225 271989
rect 64259 271961 64287 271989
rect 64321 271961 64349 271989
rect 64383 271961 64411 271989
rect 66057 299058 66085 299086
rect 66119 299058 66147 299086
rect 66181 299058 66209 299086
rect 66243 299058 66271 299086
rect 66057 298996 66085 299024
rect 66119 298996 66147 299024
rect 66181 298996 66209 299024
rect 66243 298996 66271 299024
rect 66057 298934 66085 298962
rect 66119 298934 66147 298962
rect 66181 298934 66209 298962
rect 66243 298934 66271 298962
rect 66057 298872 66085 298900
rect 66119 298872 66147 298900
rect 66181 298872 66209 298900
rect 66243 298872 66271 298900
rect 66057 293147 66085 293175
rect 66119 293147 66147 293175
rect 66181 293147 66209 293175
rect 66243 293147 66271 293175
rect 66057 293085 66085 293113
rect 66119 293085 66147 293113
rect 66181 293085 66209 293113
rect 66243 293085 66271 293113
rect 66057 293023 66085 293051
rect 66119 293023 66147 293051
rect 66181 293023 66209 293051
rect 66243 293023 66271 293051
rect 66057 292961 66085 292989
rect 66119 292961 66147 292989
rect 66181 292961 66209 292989
rect 66243 292961 66271 292989
rect 66057 284147 66085 284175
rect 66119 284147 66147 284175
rect 66181 284147 66209 284175
rect 66243 284147 66271 284175
rect 66057 284085 66085 284113
rect 66119 284085 66147 284113
rect 66181 284085 66209 284113
rect 66243 284085 66271 284113
rect 66057 284023 66085 284051
rect 66119 284023 66147 284051
rect 66181 284023 66209 284051
rect 66243 284023 66271 284051
rect 66057 283961 66085 283989
rect 66119 283961 66147 283989
rect 66181 283961 66209 283989
rect 66243 283961 66271 283989
rect 66057 275147 66085 275175
rect 66119 275147 66147 275175
rect 66181 275147 66209 275175
rect 66243 275147 66271 275175
rect 66057 275085 66085 275113
rect 66119 275085 66147 275113
rect 66181 275085 66209 275113
rect 66243 275085 66271 275113
rect 66057 275023 66085 275051
rect 66119 275023 66147 275051
rect 66181 275023 66209 275051
rect 66243 275023 66271 275051
rect 66057 274961 66085 274989
rect 66119 274961 66147 274989
rect 66181 274961 66209 274989
rect 66243 274961 66271 274989
rect 79557 298578 79585 298606
rect 79619 298578 79647 298606
rect 79681 298578 79709 298606
rect 79743 298578 79771 298606
rect 79557 298516 79585 298544
rect 79619 298516 79647 298544
rect 79681 298516 79709 298544
rect 79743 298516 79771 298544
rect 79557 298454 79585 298482
rect 79619 298454 79647 298482
rect 79681 298454 79709 298482
rect 79743 298454 79771 298482
rect 79557 298392 79585 298420
rect 79619 298392 79647 298420
rect 79681 298392 79709 298420
rect 79743 298392 79771 298420
rect 79557 290147 79585 290175
rect 79619 290147 79647 290175
rect 79681 290147 79709 290175
rect 79743 290147 79771 290175
rect 79557 290085 79585 290113
rect 79619 290085 79647 290113
rect 79681 290085 79709 290113
rect 79743 290085 79771 290113
rect 79557 290023 79585 290051
rect 79619 290023 79647 290051
rect 79681 290023 79709 290051
rect 79743 290023 79771 290051
rect 79557 289961 79585 289989
rect 79619 289961 79647 289989
rect 79681 289961 79709 289989
rect 79743 289961 79771 289989
rect 79557 281147 79585 281175
rect 79619 281147 79647 281175
rect 79681 281147 79709 281175
rect 79743 281147 79771 281175
rect 79557 281085 79585 281113
rect 79619 281085 79647 281113
rect 79681 281085 79709 281113
rect 79743 281085 79771 281113
rect 79557 281023 79585 281051
rect 79619 281023 79647 281051
rect 79681 281023 79709 281051
rect 79743 281023 79771 281051
rect 79557 280961 79585 280989
rect 79619 280961 79647 280989
rect 79681 280961 79709 280989
rect 79743 280961 79771 280989
rect 79557 272147 79585 272175
rect 79619 272147 79647 272175
rect 79681 272147 79709 272175
rect 79743 272147 79771 272175
rect 79557 272085 79585 272113
rect 79619 272085 79647 272113
rect 79681 272085 79709 272113
rect 79743 272085 79771 272113
rect 79557 272023 79585 272051
rect 79619 272023 79647 272051
rect 79681 272023 79709 272051
rect 79743 272023 79771 272051
rect 79557 271961 79585 271989
rect 79619 271961 79647 271989
rect 79681 271961 79709 271989
rect 79743 271961 79771 271989
rect 81417 299058 81445 299086
rect 81479 299058 81507 299086
rect 81541 299058 81569 299086
rect 81603 299058 81631 299086
rect 81417 298996 81445 299024
rect 81479 298996 81507 299024
rect 81541 298996 81569 299024
rect 81603 298996 81631 299024
rect 81417 298934 81445 298962
rect 81479 298934 81507 298962
rect 81541 298934 81569 298962
rect 81603 298934 81631 298962
rect 81417 298872 81445 298900
rect 81479 298872 81507 298900
rect 81541 298872 81569 298900
rect 81603 298872 81631 298900
rect 81417 293147 81445 293175
rect 81479 293147 81507 293175
rect 81541 293147 81569 293175
rect 81603 293147 81631 293175
rect 81417 293085 81445 293113
rect 81479 293085 81507 293113
rect 81541 293085 81569 293113
rect 81603 293085 81631 293113
rect 81417 293023 81445 293051
rect 81479 293023 81507 293051
rect 81541 293023 81569 293051
rect 81603 293023 81631 293051
rect 81417 292961 81445 292989
rect 81479 292961 81507 292989
rect 81541 292961 81569 292989
rect 81603 292961 81631 292989
rect 81417 284147 81445 284175
rect 81479 284147 81507 284175
rect 81541 284147 81569 284175
rect 81603 284147 81631 284175
rect 81417 284085 81445 284113
rect 81479 284085 81507 284113
rect 81541 284085 81569 284113
rect 81603 284085 81631 284113
rect 81417 284023 81445 284051
rect 81479 284023 81507 284051
rect 81541 284023 81569 284051
rect 81603 284023 81631 284051
rect 81417 283961 81445 283989
rect 81479 283961 81507 283989
rect 81541 283961 81569 283989
rect 81603 283961 81631 283989
rect 81417 275147 81445 275175
rect 81479 275147 81507 275175
rect 81541 275147 81569 275175
rect 81603 275147 81631 275175
rect 81417 275085 81445 275113
rect 81479 275085 81507 275113
rect 81541 275085 81569 275113
rect 81603 275085 81631 275113
rect 81417 275023 81445 275051
rect 81479 275023 81507 275051
rect 81541 275023 81569 275051
rect 81603 275023 81631 275051
rect 81417 274961 81445 274989
rect 81479 274961 81507 274989
rect 81541 274961 81569 274989
rect 81603 274961 81631 274989
rect 94917 298578 94945 298606
rect 94979 298578 95007 298606
rect 95041 298578 95069 298606
rect 95103 298578 95131 298606
rect 94917 298516 94945 298544
rect 94979 298516 95007 298544
rect 95041 298516 95069 298544
rect 95103 298516 95131 298544
rect 94917 298454 94945 298482
rect 94979 298454 95007 298482
rect 95041 298454 95069 298482
rect 95103 298454 95131 298482
rect 94917 298392 94945 298420
rect 94979 298392 95007 298420
rect 95041 298392 95069 298420
rect 95103 298392 95131 298420
rect 94917 290147 94945 290175
rect 94979 290147 95007 290175
rect 95041 290147 95069 290175
rect 95103 290147 95131 290175
rect 94917 290085 94945 290113
rect 94979 290085 95007 290113
rect 95041 290085 95069 290113
rect 95103 290085 95131 290113
rect 94917 290023 94945 290051
rect 94979 290023 95007 290051
rect 95041 290023 95069 290051
rect 95103 290023 95131 290051
rect 94917 289961 94945 289989
rect 94979 289961 95007 289989
rect 95041 289961 95069 289989
rect 95103 289961 95131 289989
rect 94917 281147 94945 281175
rect 94979 281147 95007 281175
rect 95041 281147 95069 281175
rect 95103 281147 95131 281175
rect 94917 281085 94945 281113
rect 94979 281085 95007 281113
rect 95041 281085 95069 281113
rect 95103 281085 95131 281113
rect 94917 281023 94945 281051
rect 94979 281023 95007 281051
rect 95041 281023 95069 281051
rect 95103 281023 95131 281051
rect 94917 280961 94945 280989
rect 94979 280961 95007 280989
rect 95041 280961 95069 280989
rect 95103 280961 95131 280989
rect 94917 272147 94945 272175
rect 94979 272147 95007 272175
rect 95041 272147 95069 272175
rect 95103 272147 95131 272175
rect 94917 272085 94945 272113
rect 94979 272085 95007 272113
rect 95041 272085 95069 272113
rect 95103 272085 95131 272113
rect 94917 272023 94945 272051
rect 94979 272023 95007 272051
rect 95041 272023 95069 272051
rect 95103 272023 95131 272051
rect 94917 271961 94945 271989
rect 94979 271961 95007 271989
rect 95041 271961 95069 271989
rect 95103 271961 95131 271989
rect 29939 266147 29967 266175
rect 30001 266147 30029 266175
rect 29939 266085 29967 266113
rect 30001 266085 30029 266113
rect 29939 266023 29967 266051
rect 30001 266023 30029 266051
rect 29939 265961 29967 265989
rect 30001 265961 30029 265989
rect 45299 266147 45327 266175
rect 45361 266147 45389 266175
rect 45299 266085 45327 266113
rect 45361 266085 45389 266113
rect 45299 266023 45327 266051
rect 45361 266023 45389 266051
rect 45299 265961 45327 265989
rect 45361 265961 45389 265989
rect 60659 266147 60687 266175
rect 60721 266147 60749 266175
rect 60659 266085 60687 266113
rect 60721 266085 60749 266113
rect 60659 266023 60687 266051
rect 60721 266023 60749 266051
rect 60659 265961 60687 265989
rect 60721 265961 60749 265989
rect 76019 266147 76047 266175
rect 76081 266147 76109 266175
rect 76019 266085 76047 266113
rect 76081 266085 76109 266113
rect 76019 266023 76047 266051
rect 76081 266023 76109 266051
rect 76019 265961 76047 265989
rect 76081 265961 76109 265989
rect 18117 263147 18145 263175
rect 18179 263147 18207 263175
rect 18241 263147 18269 263175
rect 18303 263147 18331 263175
rect 18117 263085 18145 263113
rect 18179 263085 18207 263113
rect 18241 263085 18269 263113
rect 18303 263085 18331 263113
rect 18117 263023 18145 263051
rect 18179 263023 18207 263051
rect 18241 263023 18269 263051
rect 18303 263023 18331 263051
rect 18117 262961 18145 262989
rect 18179 262961 18207 262989
rect 18241 262961 18269 262989
rect 18303 262961 18331 262989
rect 22259 263147 22287 263175
rect 22321 263147 22349 263175
rect 22259 263085 22287 263113
rect 22321 263085 22349 263113
rect 22259 263023 22287 263051
rect 22321 263023 22349 263051
rect 22259 262961 22287 262989
rect 22321 262961 22349 262989
rect 37619 263147 37647 263175
rect 37681 263147 37709 263175
rect 37619 263085 37647 263113
rect 37681 263085 37709 263113
rect 37619 263023 37647 263051
rect 37681 263023 37709 263051
rect 37619 262961 37647 262989
rect 37681 262961 37709 262989
rect 52979 263147 53007 263175
rect 53041 263147 53069 263175
rect 52979 263085 53007 263113
rect 53041 263085 53069 263113
rect 52979 263023 53007 263051
rect 53041 263023 53069 263051
rect 52979 262961 53007 262989
rect 53041 262961 53069 262989
rect 68339 263147 68367 263175
rect 68401 263147 68429 263175
rect 68339 263085 68367 263113
rect 68401 263085 68429 263113
rect 68339 263023 68367 263051
rect 68401 263023 68429 263051
rect 68339 262961 68367 262989
rect 68401 262961 68429 262989
rect 83699 263147 83727 263175
rect 83761 263147 83789 263175
rect 83699 263085 83727 263113
rect 83761 263085 83789 263113
rect 83699 263023 83727 263051
rect 83761 263023 83789 263051
rect 83699 262961 83727 262989
rect 83761 262961 83789 262989
rect 94917 263147 94945 263175
rect 94979 263147 95007 263175
rect 95041 263147 95069 263175
rect 95103 263147 95131 263175
rect 94917 263085 94945 263113
rect 94979 263085 95007 263113
rect 95041 263085 95069 263113
rect 95103 263085 95131 263113
rect 94917 263023 94945 263051
rect 94979 263023 95007 263051
rect 95041 263023 95069 263051
rect 95103 263023 95131 263051
rect 94917 262961 94945 262989
rect 94979 262961 95007 262989
rect 95041 262961 95069 262989
rect 95103 262961 95131 262989
rect 29939 257147 29967 257175
rect 30001 257147 30029 257175
rect 29939 257085 29967 257113
rect 30001 257085 30029 257113
rect 29939 257023 29967 257051
rect 30001 257023 30029 257051
rect 29939 256961 29967 256989
rect 30001 256961 30029 256989
rect 45299 257147 45327 257175
rect 45361 257147 45389 257175
rect 45299 257085 45327 257113
rect 45361 257085 45389 257113
rect 45299 257023 45327 257051
rect 45361 257023 45389 257051
rect 45299 256961 45327 256989
rect 45361 256961 45389 256989
rect 60659 257147 60687 257175
rect 60721 257147 60749 257175
rect 60659 257085 60687 257113
rect 60721 257085 60749 257113
rect 60659 257023 60687 257051
rect 60721 257023 60749 257051
rect 60659 256961 60687 256989
rect 60721 256961 60749 256989
rect 76019 257147 76047 257175
rect 76081 257147 76109 257175
rect 76019 257085 76047 257113
rect 76081 257085 76109 257113
rect 76019 257023 76047 257051
rect 76081 257023 76109 257051
rect 76019 256961 76047 256989
rect 76081 256961 76109 256989
rect 18117 254147 18145 254175
rect 18179 254147 18207 254175
rect 18241 254147 18269 254175
rect 18303 254147 18331 254175
rect 18117 254085 18145 254113
rect 18179 254085 18207 254113
rect 18241 254085 18269 254113
rect 18303 254085 18331 254113
rect 18117 254023 18145 254051
rect 18179 254023 18207 254051
rect 18241 254023 18269 254051
rect 18303 254023 18331 254051
rect 18117 253961 18145 253989
rect 18179 253961 18207 253989
rect 18241 253961 18269 253989
rect 18303 253961 18331 253989
rect 22259 254147 22287 254175
rect 22321 254147 22349 254175
rect 22259 254085 22287 254113
rect 22321 254085 22349 254113
rect 22259 254023 22287 254051
rect 22321 254023 22349 254051
rect 22259 253961 22287 253989
rect 22321 253961 22349 253989
rect 37619 254147 37647 254175
rect 37681 254147 37709 254175
rect 37619 254085 37647 254113
rect 37681 254085 37709 254113
rect 37619 254023 37647 254051
rect 37681 254023 37709 254051
rect 37619 253961 37647 253989
rect 37681 253961 37709 253989
rect 52979 254147 53007 254175
rect 53041 254147 53069 254175
rect 52979 254085 53007 254113
rect 53041 254085 53069 254113
rect 52979 254023 53007 254051
rect 53041 254023 53069 254051
rect 52979 253961 53007 253989
rect 53041 253961 53069 253989
rect 68339 254147 68367 254175
rect 68401 254147 68429 254175
rect 68339 254085 68367 254113
rect 68401 254085 68429 254113
rect 68339 254023 68367 254051
rect 68401 254023 68429 254051
rect 68339 253961 68367 253989
rect 68401 253961 68429 253989
rect 83699 254147 83727 254175
rect 83761 254147 83789 254175
rect 83699 254085 83727 254113
rect 83761 254085 83789 254113
rect 83699 254023 83727 254051
rect 83761 254023 83789 254051
rect 83699 253961 83727 253989
rect 83761 253961 83789 253989
rect 94917 254147 94945 254175
rect 94979 254147 95007 254175
rect 95041 254147 95069 254175
rect 95103 254147 95131 254175
rect 94917 254085 94945 254113
rect 94979 254085 95007 254113
rect 95041 254085 95069 254113
rect 95103 254085 95131 254113
rect 94917 254023 94945 254051
rect 94979 254023 95007 254051
rect 95041 254023 95069 254051
rect 95103 254023 95131 254051
rect 94917 253961 94945 253989
rect 94979 253961 95007 253989
rect 95041 253961 95069 253989
rect 95103 253961 95131 253989
rect 29939 248147 29967 248175
rect 30001 248147 30029 248175
rect 29939 248085 29967 248113
rect 30001 248085 30029 248113
rect 29939 248023 29967 248051
rect 30001 248023 30029 248051
rect 29939 247961 29967 247989
rect 30001 247961 30029 247989
rect 45299 248147 45327 248175
rect 45361 248147 45389 248175
rect 45299 248085 45327 248113
rect 45361 248085 45389 248113
rect 45299 248023 45327 248051
rect 45361 248023 45389 248051
rect 45299 247961 45327 247989
rect 45361 247961 45389 247989
rect 60659 248147 60687 248175
rect 60721 248147 60749 248175
rect 60659 248085 60687 248113
rect 60721 248085 60749 248113
rect 60659 248023 60687 248051
rect 60721 248023 60749 248051
rect 60659 247961 60687 247989
rect 60721 247961 60749 247989
rect 76019 248147 76047 248175
rect 76081 248147 76109 248175
rect 76019 248085 76047 248113
rect 76081 248085 76109 248113
rect 76019 248023 76047 248051
rect 76081 248023 76109 248051
rect 76019 247961 76047 247989
rect 76081 247961 76109 247989
rect 18117 245147 18145 245175
rect 18179 245147 18207 245175
rect 18241 245147 18269 245175
rect 18303 245147 18331 245175
rect 18117 245085 18145 245113
rect 18179 245085 18207 245113
rect 18241 245085 18269 245113
rect 18303 245085 18331 245113
rect 18117 245023 18145 245051
rect 18179 245023 18207 245051
rect 18241 245023 18269 245051
rect 18303 245023 18331 245051
rect 18117 244961 18145 244989
rect 18179 244961 18207 244989
rect 18241 244961 18269 244989
rect 18303 244961 18331 244989
rect 22259 245147 22287 245175
rect 22321 245147 22349 245175
rect 22259 245085 22287 245113
rect 22321 245085 22349 245113
rect 22259 245023 22287 245051
rect 22321 245023 22349 245051
rect 22259 244961 22287 244989
rect 22321 244961 22349 244989
rect 37619 245147 37647 245175
rect 37681 245147 37709 245175
rect 37619 245085 37647 245113
rect 37681 245085 37709 245113
rect 37619 245023 37647 245051
rect 37681 245023 37709 245051
rect 37619 244961 37647 244989
rect 37681 244961 37709 244989
rect 52979 245147 53007 245175
rect 53041 245147 53069 245175
rect 52979 245085 53007 245113
rect 53041 245085 53069 245113
rect 52979 245023 53007 245051
rect 53041 245023 53069 245051
rect 52979 244961 53007 244989
rect 53041 244961 53069 244989
rect 68339 245147 68367 245175
rect 68401 245147 68429 245175
rect 68339 245085 68367 245113
rect 68401 245085 68429 245113
rect 68339 245023 68367 245051
rect 68401 245023 68429 245051
rect 68339 244961 68367 244989
rect 68401 244961 68429 244989
rect 83699 245147 83727 245175
rect 83761 245147 83789 245175
rect 83699 245085 83727 245113
rect 83761 245085 83789 245113
rect 83699 245023 83727 245051
rect 83761 245023 83789 245051
rect 83699 244961 83727 244989
rect 83761 244961 83789 244989
rect 94917 245147 94945 245175
rect 94979 245147 95007 245175
rect 95041 245147 95069 245175
rect 95103 245147 95131 245175
rect 94917 245085 94945 245113
rect 94979 245085 95007 245113
rect 95041 245085 95069 245113
rect 95103 245085 95131 245113
rect 94917 245023 94945 245051
rect 94979 245023 95007 245051
rect 95041 245023 95069 245051
rect 95103 245023 95131 245051
rect 94917 244961 94945 244989
rect 94979 244961 95007 244989
rect 95041 244961 95069 244989
rect 95103 244961 95131 244989
rect 29939 239147 29967 239175
rect 30001 239147 30029 239175
rect 29939 239085 29967 239113
rect 30001 239085 30029 239113
rect 29939 239023 29967 239051
rect 30001 239023 30029 239051
rect 29939 238961 29967 238989
rect 30001 238961 30029 238989
rect 45299 239147 45327 239175
rect 45361 239147 45389 239175
rect 45299 239085 45327 239113
rect 45361 239085 45389 239113
rect 45299 239023 45327 239051
rect 45361 239023 45389 239051
rect 45299 238961 45327 238989
rect 45361 238961 45389 238989
rect 60659 239147 60687 239175
rect 60721 239147 60749 239175
rect 60659 239085 60687 239113
rect 60721 239085 60749 239113
rect 60659 239023 60687 239051
rect 60721 239023 60749 239051
rect 60659 238961 60687 238989
rect 60721 238961 60749 238989
rect 76019 239147 76047 239175
rect 76081 239147 76109 239175
rect 76019 239085 76047 239113
rect 76081 239085 76109 239113
rect 76019 239023 76047 239051
rect 76081 239023 76109 239051
rect 76019 238961 76047 238989
rect 76081 238961 76109 238989
rect 18117 236147 18145 236175
rect 18179 236147 18207 236175
rect 18241 236147 18269 236175
rect 18303 236147 18331 236175
rect 18117 236085 18145 236113
rect 18179 236085 18207 236113
rect 18241 236085 18269 236113
rect 18303 236085 18331 236113
rect 18117 236023 18145 236051
rect 18179 236023 18207 236051
rect 18241 236023 18269 236051
rect 18303 236023 18331 236051
rect 18117 235961 18145 235989
rect 18179 235961 18207 235989
rect 18241 235961 18269 235989
rect 18303 235961 18331 235989
rect 22259 236147 22287 236175
rect 22321 236147 22349 236175
rect 22259 236085 22287 236113
rect 22321 236085 22349 236113
rect 22259 236023 22287 236051
rect 22321 236023 22349 236051
rect 22259 235961 22287 235989
rect 22321 235961 22349 235989
rect 37619 236147 37647 236175
rect 37681 236147 37709 236175
rect 37619 236085 37647 236113
rect 37681 236085 37709 236113
rect 37619 236023 37647 236051
rect 37681 236023 37709 236051
rect 37619 235961 37647 235989
rect 37681 235961 37709 235989
rect 52979 236147 53007 236175
rect 53041 236147 53069 236175
rect 52979 236085 53007 236113
rect 53041 236085 53069 236113
rect 52979 236023 53007 236051
rect 53041 236023 53069 236051
rect 52979 235961 53007 235989
rect 53041 235961 53069 235989
rect 68339 236147 68367 236175
rect 68401 236147 68429 236175
rect 68339 236085 68367 236113
rect 68401 236085 68429 236113
rect 68339 236023 68367 236051
rect 68401 236023 68429 236051
rect 68339 235961 68367 235989
rect 68401 235961 68429 235989
rect 83699 236147 83727 236175
rect 83761 236147 83789 236175
rect 83699 236085 83727 236113
rect 83761 236085 83789 236113
rect 83699 236023 83727 236051
rect 83761 236023 83789 236051
rect 83699 235961 83727 235989
rect 83761 235961 83789 235989
rect 94917 236147 94945 236175
rect 94979 236147 95007 236175
rect 95041 236147 95069 236175
rect 95103 236147 95131 236175
rect 94917 236085 94945 236113
rect 94979 236085 95007 236113
rect 95041 236085 95069 236113
rect 95103 236085 95131 236113
rect 94917 236023 94945 236051
rect 94979 236023 95007 236051
rect 95041 236023 95069 236051
rect 95103 236023 95131 236051
rect 94917 235961 94945 235989
rect 94979 235961 95007 235989
rect 95041 235961 95069 235989
rect 95103 235961 95131 235989
rect 29939 230147 29967 230175
rect 30001 230147 30029 230175
rect 29939 230085 29967 230113
rect 30001 230085 30029 230113
rect 29939 230023 29967 230051
rect 30001 230023 30029 230051
rect 29939 229961 29967 229989
rect 30001 229961 30029 229989
rect 45299 230147 45327 230175
rect 45361 230147 45389 230175
rect 45299 230085 45327 230113
rect 45361 230085 45389 230113
rect 45299 230023 45327 230051
rect 45361 230023 45389 230051
rect 45299 229961 45327 229989
rect 45361 229961 45389 229989
rect 60659 230147 60687 230175
rect 60721 230147 60749 230175
rect 60659 230085 60687 230113
rect 60721 230085 60749 230113
rect 60659 230023 60687 230051
rect 60721 230023 60749 230051
rect 60659 229961 60687 229989
rect 60721 229961 60749 229989
rect 76019 230147 76047 230175
rect 76081 230147 76109 230175
rect 76019 230085 76047 230113
rect 76081 230085 76109 230113
rect 76019 230023 76047 230051
rect 76081 230023 76109 230051
rect 76019 229961 76047 229989
rect 76081 229961 76109 229989
rect 18117 227147 18145 227175
rect 18179 227147 18207 227175
rect 18241 227147 18269 227175
rect 18303 227147 18331 227175
rect 18117 227085 18145 227113
rect 18179 227085 18207 227113
rect 18241 227085 18269 227113
rect 18303 227085 18331 227113
rect 18117 227023 18145 227051
rect 18179 227023 18207 227051
rect 18241 227023 18269 227051
rect 18303 227023 18331 227051
rect 18117 226961 18145 226989
rect 18179 226961 18207 226989
rect 18241 226961 18269 226989
rect 18303 226961 18331 226989
rect 22259 227147 22287 227175
rect 22321 227147 22349 227175
rect 22259 227085 22287 227113
rect 22321 227085 22349 227113
rect 22259 227023 22287 227051
rect 22321 227023 22349 227051
rect 22259 226961 22287 226989
rect 22321 226961 22349 226989
rect 37619 227147 37647 227175
rect 37681 227147 37709 227175
rect 37619 227085 37647 227113
rect 37681 227085 37709 227113
rect 37619 227023 37647 227051
rect 37681 227023 37709 227051
rect 37619 226961 37647 226989
rect 37681 226961 37709 226989
rect 52979 227147 53007 227175
rect 53041 227147 53069 227175
rect 52979 227085 53007 227113
rect 53041 227085 53069 227113
rect 52979 227023 53007 227051
rect 53041 227023 53069 227051
rect 52979 226961 53007 226989
rect 53041 226961 53069 226989
rect 68339 227147 68367 227175
rect 68401 227147 68429 227175
rect 68339 227085 68367 227113
rect 68401 227085 68429 227113
rect 68339 227023 68367 227051
rect 68401 227023 68429 227051
rect 68339 226961 68367 226989
rect 68401 226961 68429 226989
rect 83699 227147 83727 227175
rect 83761 227147 83789 227175
rect 83699 227085 83727 227113
rect 83761 227085 83789 227113
rect 83699 227023 83727 227051
rect 83761 227023 83789 227051
rect 83699 226961 83727 226989
rect 83761 226961 83789 226989
rect 94917 227147 94945 227175
rect 94979 227147 95007 227175
rect 95041 227147 95069 227175
rect 95103 227147 95131 227175
rect 94917 227085 94945 227113
rect 94979 227085 95007 227113
rect 95041 227085 95069 227113
rect 95103 227085 95131 227113
rect 94917 227023 94945 227051
rect 94979 227023 95007 227051
rect 95041 227023 95069 227051
rect 95103 227023 95131 227051
rect 94917 226961 94945 226989
rect 94979 226961 95007 226989
rect 95041 226961 95069 226989
rect 95103 226961 95131 226989
rect 29939 221147 29967 221175
rect 30001 221147 30029 221175
rect 29939 221085 29967 221113
rect 30001 221085 30029 221113
rect 29939 221023 29967 221051
rect 30001 221023 30029 221051
rect 29939 220961 29967 220989
rect 30001 220961 30029 220989
rect 45299 221147 45327 221175
rect 45361 221147 45389 221175
rect 45299 221085 45327 221113
rect 45361 221085 45389 221113
rect 45299 221023 45327 221051
rect 45361 221023 45389 221051
rect 45299 220961 45327 220989
rect 45361 220961 45389 220989
rect 60659 221147 60687 221175
rect 60721 221147 60749 221175
rect 60659 221085 60687 221113
rect 60721 221085 60749 221113
rect 60659 221023 60687 221051
rect 60721 221023 60749 221051
rect 60659 220961 60687 220989
rect 60721 220961 60749 220989
rect 76019 221147 76047 221175
rect 76081 221147 76109 221175
rect 76019 221085 76047 221113
rect 76081 221085 76109 221113
rect 76019 221023 76047 221051
rect 76081 221023 76109 221051
rect 76019 220961 76047 220989
rect 76081 220961 76109 220989
rect 18117 218147 18145 218175
rect 18179 218147 18207 218175
rect 18241 218147 18269 218175
rect 18303 218147 18331 218175
rect 18117 218085 18145 218113
rect 18179 218085 18207 218113
rect 18241 218085 18269 218113
rect 18303 218085 18331 218113
rect 18117 218023 18145 218051
rect 18179 218023 18207 218051
rect 18241 218023 18269 218051
rect 18303 218023 18331 218051
rect 18117 217961 18145 217989
rect 18179 217961 18207 217989
rect 18241 217961 18269 217989
rect 18303 217961 18331 217989
rect 22259 218147 22287 218175
rect 22321 218147 22349 218175
rect 22259 218085 22287 218113
rect 22321 218085 22349 218113
rect 22259 218023 22287 218051
rect 22321 218023 22349 218051
rect 22259 217961 22287 217989
rect 22321 217961 22349 217989
rect 37619 218147 37647 218175
rect 37681 218147 37709 218175
rect 37619 218085 37647 218113
rect 37681 218085 37709 218113
rect 37619 218023 37647 218051
rect 37681 218023 37709 218051
rect 37619 217961 37647 217989
rect 37681 217961 37709 217989
rect 52979 218147 53007 218175
rect 53041 218147 53069 218175
rect 52979 218085 53007 218113
rect 53041 218085 53069 218113
rect 52979 218023 53007 218051
rect 53041 218023 53069 218051
rect 52979 217961 53007 217989
rect 53041 217961 53069 217989
rect 68339 218147 68367 218175
rect 68401 218147 68429 218175
rect 68339 218085 68367 218113
rect 68401 218085 68429 218113
rect 68339 218023 68367 218051
rect 68401 218023 68429 218051
rect 68339 217961 68367 217989
rect 68401 217961 68429 217989
rect 83699 218147 83727 218175
rect 83761 218147 83789 218175
rect 83699 218085 83727 218113
rect 83761 218085 83789 218113
rect 83699 218023 83727 218051
rect 83761 218023 83789 218051
rect 83699 217961 83727 217989
rect 83761 217961 83789 217989
rect 94917 218147 94945 218175
rect 94979 218147 95007 218175
rect 95041 218147 95069 218175
rect 95103 218147 95131 218175
rect 94917 218085 94945 218113
rect 94979 218085 95007 218113
rect 95041 218085 95069 218113
rect 95103 218085 95131 218113
rect 94917 218023 94945 218051
rect 94979 218023 95007 218051
rect 95041 218023 95069 218051
rect 95103 218023 95131 218051
rect 94917 217961 94945 217989
rect 94979 217961 95007 217989
rect 95041 217961 95069 217989
rect 95103 217961 95131 217989
rect 29939 212147 29967 212175
rect 30001 212147 30029 212175
rect 29939 212085 29967 212113
rect 30001 212085 30029 212113
rect 29939 212023 29967 212051
rect 30001 212023 30029 212051
rect 29939 211961 29967 211989
rect 30001 211961 30029 211989
rect 45299 212147 45327 212175
rect 45361 212147 45389 212175
rect 45299 212085 45327 212113
rect 45361 212085 45389 212113
rect 45299 212023 45327 212051
rect 45361 212023 45389 212051
rect 45299 211961 45327 211989
rect 45361 211961 45389 211989
rect 60659 212147 60687 212175
rect 60721 212147 60749 212175
rect 60659 212085 60687 212113
rect 60721 212085 60749 212113
rect 60659 212023 60687 212051
rect 60721 212023 60749 212051
rect 60659 211961 60687 211989
rect 60721 211961 60749 211989
rect 76019 212147 76047 212175
rect 76081 212147 76109 212175
rect 76019 212085 76047 212113
rect 76081 212085 76109 212113
rect 76019 212023 76047 212051
rect 76081 212023 76109 212051
rect 76019 211961 76047 211989
rect 76081 211961 76109 211989
rect 18117 209147 18145 209175
rect 18179 209147 18207 209175
rect 18241 209147 18269 209175
rect 18303 209147 18331 209175
rect 18117 209085 18145 209113
rect 18179 209085 18207 209113
rect 18241 209085 18269 209113
rect 18303 209085 18331 209113
rect 18117 209023 18145 209051
rect 18179 209023 18207 209051
rect 18241 209023 18269 209051
rect 18303 209023 18331 209051
rect 18117 208961 18145 208989
rect 18179 208961 18207 208989
rect 18241 208961 18269 208989
rect 18303 208961 18331 208989
rect 22259 209147 22287 209175
rect 22321 209147 22349 209175
rect 22259 209085 22287 209113
rect 22321 209085 22349 209113
rect 22259 209023 22287 209051
rect 22321 209023 22349 209051
rect 22259 208961 22287 208989
rect 22321 208961 22349 208989
rect 37619 209147 37647 209175
rect 37681 209147 37709 209175
rect 37619 209085 37647 209113
rect 37681 209085 37709 209113
rect 37619 209023 37647 209051
rect 37681 209023 37709 209051
rect 37619 208961 37647 208989
rect 37681 208961 37709 208989
rect 52979 209147 53007 209175
rect 53041 209147 53069 209175
rect 52979 209085 53007 209113
rect 53041 209085 53069 209113
rect 52979 209023 53007 209051
rect 53041 209023 53069 209051
rect 52979 208961 53007 208989
rect 53041 208961 53069 208989
rect 68339 209147 68367 209175
rect 68401 209147 68429 209175
rect 68339 209085 68367 209113
rect 68401 209085 68429 209113
rect 68339 209023 68367 209051
rect 68401 209023 68429 209051
rect 68339 208961 68367 208989
rect 68401 208961 68429 208989
rect 83699 209147 83727 209175
rect 83761 209147 83789 209175
rect 83699 209085 83727 209113
rect 83761 209085 83789 209113
rect 83699 209023 83727 209051
rect 83761 209023 83789 209051
rect 83699 208961 83727 208989
rect 83761 208961 83789 208989
rect 94917 209147 94945 209175
rect 94979 209147 95007 209175
rect 95041 209147 95069 209175
rect 95103 209147 95131 209175
rect 94917 209085 94945 209113
rect 94979 209085 95007 209113
rect 95041 209085 95069 209113
rect 95103 209085 95131 209113
rect 94917 209023 94945 209051
rect 94979 209023 95007 209051
rect 95041 209023 95069 209051
rect 95103 209023 95131 209051
rect 94917 208961 94945 208989
rect 94979 208961 95007 208989
rect 95041 208961 95069 208989
rect 95103 208961 95131 208989
rect 29939 203147 29967 203175
rect 30001 203147 30029 203175
rect 29939 203085 29967 203113
rect 30001 203085 30029 203113
rect 29939 203023 29967 203051
rect 30001 203023 30029 203051
rect 29939 202961 29967 202989
rect 30001 202961 30029 202989
rect 45299 203147 45327 203175
rect 45361 203147 45389 203175
rect 45299 203085 45327 203113
rect 45361 203085 45389 203113
rect 45299 203023 45327 203051
rect 45361 203023 45389 203051
rect 45299 202961 45327 202989
rect 45361 202961 45389 202989
rect 60659 203147 60687 203175
rect 60721 203147 60749 203175
rect 60659 203085 60687 203113
rect 60721 203085 60749 203113
rect 60659 203023 60687 203051
rect 60721 203023 60749 203051
rect 60659 202961 60687 202989
rect 60721 202961 60749 202989
rect 76019 203147 76047 203175
rect 76081 203147 76109 203175
rect 76019 203085 76047 203113
rect 76081 203085 76109 203113
rect 76019 203023 76047 203051
rect 76081 203023 76109 203051
rect 76019 202961 76047 202989
rect 76081 202961 76109 202989
rect 18117 200147 18145 200175
rect 18179 200147 18207 200175
rect 18241 200147 18269 200175
rect 18303 200147 18331 200175
rect 18117 200085 18145 200113
rect 18179 200085 18207 200113
rect 18241 200085 18269 200113
rect 18303 200085 18331 200113
rect 18117 200023 18145 200051
rect 18179 200023 18207 200051
rect 18241 200023 18269 200051
rect 18303 200023 18331 200051
rect 18117 199961 18145 199989
rect 18179 199961 18207 199989
rect 18241 199961 18269 199989
rect 18303 199961 18331 199989
rect 22259 200147 22287 200175
rect 22321 200147 22349 200175
rect 22259 200085 22287 200113
rect 22321 200085 22349 200113
rect 22259 200023 22287 200051
rect 22321 200023 22349 200051
rect 22259 199961 22287 199989
rect 22321 199961 22349 199989
rect 37619 200147 37647 200175
rect 37681 200147 37709 200175
rect 37619 200085 37647 200113
rect 37681 200085 37709 200113
rect 37619 200023 37647 200051
rect 37681 200023 37709 200051
rect 37619 199961 37647 199989
rect 37681 199961 37709 199989
rect 52979 200147 53007 200175
rect 53041 200147 53069 200175
rect 52979 200085 53007 200113
rect 53041 200085 53069 200113
rect 52979 200023 53007 200051
rect 53041 200023 53069 200051
rect 52979 199961 53007 199989
rect 53041 199961 53069 199989
rect 68339 200147 68367 200175
rect 68401 200147 68429 200175
rect 68339 200085 68367 200113
rect 68401 200085 68429 200113
rect 68339 200023 68367 200051
rect 68401 200023 68429 200051
rect 68339 199961 68367 199989
rect 68401 199961 68429 199989
rect 83699 200147 83727 200175
rect 83761 200147 83789 200175
rect 83699 200085 83727 200113
rect 83761 200085 83789 200113
rect 83699 200023 83727 200051
rect 83761 200023 83789 200051
rect 83699 199961 83727 199989
rect 83761 199961 83789 199989
rect 94917 200147 94945 200175
rect 94979 200147 95007 200175
rect 95041 200147 95069 200175
rect 95103 200147 95131 200175
rect 94917 200085 94945 200113
rect 94979 200085 95007 200113
rect 95041 200085 95069 200113
rect 95103 200085 95131 200113
rect 94917 200023 94945 200051
rect 94979 200023 95007 200051
rect 95041 200023 95069 200051
rect 95103 200023 95131 200051
rect 94917 199961 94945 199989
rect 94979 199961 95007 199989
rect 95041 199961 95069 199989
rect 95103 199961 95131 199989
rect 29939 194147 29967 194175
rect 30001 194147 30029 194175
rect 29939 194085 29967 194113
rect 30001 194085 30029 194113
rect 29939 194023 29967 194051
rect 30001 194023 30029 194051
rect 29939 193961 29967 193989
rect 30001 193961 30029 193989
rect 45299 194147 45327 194175
rect 45361 194147 45389 194175
rect 45299 194085 45327 194113
rect 45361 194085 45389 194113
rect 45299 194023 45327 194051
rect 45361 194023 45389 194051
rect 45299 193961 45327 193989
rect 45361 193961 45389 193989
rect 60659 194147 60687 194175
rect 60721 194147 60749 194175
rect 60659 194085 60687 194113
rect 60721 194085 60749 194113
rect 60659 194023 60687 194051
rect 60721 194023 60749 194051
rect 60659 193961 60687 193989
rect 60721 193961 60749 193989
rect 76019 194147 76047 194175
rect 76081 194147 76109 194175
rect 76019 194085 76047 194113
rect 76081 194085 76109 194113
rect 76019 194023 76047 194051
rect 76081 194023 76109 194051
rect 76019 193961 76047 193989
rect 76081 193961 76109 193989
rect 18117 191147 18145 191175
rect 18179 191147 18207 191175
rect 18241 191147 18269 191175
rect 18303 191147 18331 191175
rect 18117 191085 18145 191113
rect 18179 191085 18207 191113
rect 18241 191085 18269 191113
rect 18303 191085 18331 191113
rect 18117 191023 18145 191051
rect 18179 191023 18207 191051
rect 18241 191023 18269 191051
rect 18303 191023 18331 191051
rect 18117 190961 18145 190989
rect 18179 190961 18207 190989
rect 18241 190961 18269 190989
rect 18303 190961 18331 190989
rect 22259 191147 22287 191175
rect 22321 191147 22349 191175
rect 22259 191085 22287 191113
rect 22321 191085 22349 191113
rect 22259 191023 22287 191051
rect 22321 191023 22349 191051
rect 22259 190961 22287 190989
rect 22321 190961 22349 190989
rect 37619 191147 37647 191175
rect 37681 191147 37709 191175
rect 37619 191085 37647 191113
rect 37681 191085 37709 191113
rect 37619 191023 37647 191051
rect 37681 191023 37709 191051
rect 37619 190961 37647 190989
rect 37681 190961 37709 190989
rect 52979 191147 53007 191175
rect 53041 191147 53069 191175
rect 52979 191085 53007 191113
rect 53041 191085 53069 191113
rect 52979 191023 53007 191051
rect 53041 191023 53069 191051
rect 52979 190961 53007 190989
rect 53041 190961 53069 190989
rect 68339 191147 68367 191175
rect 68401 191147 68429 191175
rect 68339 191085 68367 191113
rect 68401 191085 68429 191113
rect 68339 191023 68367 191051
rect 68401 191023 68429 191051
rect 68339 190961 68367 190989
rect 68401 190961 68429 190989
rect 83699 191147 83727 191175
rect 83761 191147 83789 191175
rect 83699 191085 83727 191113
rect 83761 191085 83789 191113
rect 83699 191023 83727 191051
rect 83761 191023 83789 191051
rect 83699 190961 83727 190989
rect 83761 190961 83789 190989
rect 94917 191147 94945 191175
rect 94979 191147 95007 191175
rect 95041 191147 95069 191175
rect 95103 191147 95131 191175
rect 94917 191085 94945 191113
rect 94979 191085 95007 191113
rect 95041 191085 95069 191113
rect 95103 191085 95131 191113
rect 94917 191023 94945 191051
rect 94979 191023 95007 191051
rect 95041 191023 95069 191051
rect 95103 191023 95131 191051
rect 94917 190961 94945 190989
rect 94979 190961 95007 190989
rect 95041 190961 95069 190989
rect 95103 190961 95131 190989
rect 29939 185147 29967 185175
rect 30001 185147 30029 185175
rect 29939 185085 29967 185113
rect 30001 185085 30029 185113
rect 29939 185023 29967 185051
rect 30001 185023 30029 185051
rect 29939 184961 29967 184989
rect 30001 184961 30029 184989
rect 45299 185147 45327 185175
rect 45361 185147 45389 185175
rect 45299 185085 45327 185113
rect 45361 185085 45389 185113
rect 45299 185023 45327 185051
rect 45361 185023 45389 185051
rect 45299 184961 45327 184989
rect 45361 184961 45389 184989
rect 60659 185147 60687 185175
rect 60721 185147 60749 185175
rect 60659 185085 60687 185113
rect 60721 185085 60749 185113
rect 60659 185023 60687 185051
rect 60721 185023 60749 185051
rect 60659 184961 60687 184989
rect 60721 184961 60749 184989
rect 76019 185147 76047 185175
rect 76081 185147 76109 185175
rect 76019 185085 76047 185113
rect 76081 185085 76109 185113
rect 76019 185023 76047 185051
rect 76081 185023 76109 185051
rect 76019 184961 76047 184989
rect 76081 184961 76109 184989
rect 18117 182147 18145 182175
rect 18179 182147 18207 182175
rect 18241 182147 18269 182175
rect 18303 182147 18331 182175
rect 18117 182085 18145 182113
rect 18179 182085 18207 182113
rect 18241 182085 18269 182113
rect 18303 182085 18331 182113
rect 18117 182023 18145 182051
rect 18179 182023 18207 182051
rect 18241 182023 18269 182051
rect 18303 182023 18331 182051
rect 18117 181961 18145 181989
rect 18179 181961 18207 181989
rect 18241 181961 18269 181989
rect 18303 181961 18331 181989
rect 22259 182147 22287 182175
rect 22321 182147 22349 182175
rect 22259 182085 22287 182113
rect 22321 182085 22349 182113
rect 22259 182023 22287 182051
rect 22321 182023 22349 182051
rect 22259 181961 22287 181989
rect 22321 181961 22349 181989
rect 37619 182147 37647 182175
rect 37681 182147 37709 182175
rect 37619 182085 37647 182113
rect 37681 182085 37709 182113
rect 37619 182023 37647 182051
rect 37681 182023 37709 182051
rect 37619 181961 37647 181989
rect 37681 181961 37709 181989
rect 52979 182147 53007 182175
rect 53041 182147 53069 182175
rect 52979 182085 53007 182113
rect 53041 182085 53069 182113
rect 52979 182023 53007 182051
rect 53041 182023 53069 182051
rect 52979 181961 53007 181989
rect 53041 181961 53069 181989
rect 68339 182147 68367 182175
rect 68401 182147 68429 182175
rect 68339 182085 68367 182113
rect 68401 182085 68429 182113
rect 68339 182023 68367 182051
rect 68401 182023 68429 182051
rect 68339 181961 68367 181989
rect 68401 181961 68429 181989
rect 83699 182147 83727 182175
rect 83761 182147 83789 182175
rect 83699 182085 83727 182113
rect 83761 182085 83789 182113
rect 83699 182023 83727 182051
rect 83761 182023 83789 182051
rect 83699 181961 83727 181989
rect 83761 181961 83789 181989
rect 94917 182147 94945 182175
rect 94979 182147 95007 182175
rect 95041 182147 95069 182175
rect 95103 182147 95131 182175
rect 94917 182085 94945 182113
rect 94979 182085 95007 182113
rect 95041 182085 95069 182113
rect 95103 182085 95131 182113
rect 94917 182023 94945 182051
rect 94979 182023 95007 182051
rect 95041 182023 95069 182051
rect 95103 182023 95131 182051
rect 94917 181961 94945 181989
rect 94979 181961 95007 181989
rect 95041 181961 95069 181989
rect 95103 181961 95131 181989
rect 29939 176147 29967 176175
rect 30001 176147 30029 176175
rect 29939 176085 29967 176113
rect 30001 176085 30029 176113
rect 29939 176023 29967 176051
rect 30001 176023 30029 176051
rect 29939 175961 29967 175989
rect 30001 175961 30029 175989
rect 45299 176147 45327 176175
rect 45361 176147 45389 176175
rect 45299 176085 45327 176113
rect 45361 176085 45389 176113
rect 45299 176023 45327 176051
rect 45361 176023 45389 176051
rect 45299 175961 45327 175989
rect 45361 175961 45389 175989
rect 60659 176147 60687 176175
rect 60721 176147 60749 176175
rect 60659 176085 60687 176113
rect 60721 176085 60749 176113
rect 60659 176023 60687 176051
rect 60721 176023 60749 176051
rect 60659 175961 60687 175989
rect 60721 175961 60749 175989
rect 76019 176147 76047 176175
rect 76081 176147 76109 176175
rect 76019 176085 76047 176113
rect 76081 176085 76109 176113
rect 76019 176023 76047 176051
rect 76081 176023 76109 176051
rect 76019 175961 76047 175989
rect 76081 175961 76109 175989
rect 18117 173147 18145 173175
rect 18179 173147 18207 173175
rect 18241 173147 18269 173175
rect 18303 173147 18331 173175
rect 18117 173085 18145 173113
rect 18179 173085 18207 173113
rect 18241 173085 18269 173113
rect 18303 173085 18331 173113
rect 18117 173023 18145 173051
rect 18179 173023 18207 173051
rect 18241 173023 18269 173051
rect 18303 173023 18331 173051
rect 18117 172961 18145 172989
rect 18179 172961 18207 172989
rect 18241 172961 18269 172989
rect 18303 172961 18331 172989
rect 22259 173147 22287 173175
rect 22321 173147 22349 173175
rect 22259 173085 22287 173113
rect 22321 173085 22349 173113
rect 22259 173023 22287 173051
rect 22321 173023 22349 173051
rect 22259 172961 22287 172989
rect 22321 172961 22349 172989
rect 37619 173147 37647 173175
rect 37681 173147 37709 173175
rect 37619 173085 37647 173113
rect 37681 173085 37709 173113
rect 37619 173023 37647 173051
rect 37681 173023 37709 173051
rect 37619 172961 37647 172989
rect 37681 172961 37709 172989
rect 52979 173147 53007 173175
rect 53041 173147 53069 173175
rect 52979 173085 53007 173113
rect 53041 173085 53069 173113
rect 52979 173023 53007 173051
rect 53041 173023 53069 173051
rect 52979 172961 53007 172989
rect 53041 172961 53069 172989
rect 68339 173147 68367 173175
rect 68401 173147 68429 173175
rect 68339 173085 68367 173113
rect 68401 173085 68429 173113
rect 68339 173023 68367 173051
rect 68401 173023 68429 173051
rect 68339 172961 68367 172989
rect 68401 172961 68429 172989
rect 83699 173147 83727 173175
rect 83761 173147 83789 173175
rect 83699 173085 83727 173113
rect 83761 173085 83789 173113
rect 83699 173023 83727 173051
rect 83761 173023 83789 173051
rect 83699 172961 83727 172989
rect 83761 172961 83789 172989
rect 94917 173147 94945 173175
rect 94979 173147 95007 173175
rect 95041 173147 95069 173175
rect 95103 173147 95131 173175
rect 94917 173085 94945 173113
rect 94979 173085 95007 173113
rect 95041 173085 95069 173113
rect 95103 173085 95131 173113
rect 94917 173023 94945 173051
rect 94979 173023 95007 173051
rect 95041 173023 95069 173051
rect 95103 173023 95131 173051
rect 94917 172961 94945 172989
rect 94979 172961 95007 172989
rect 95041 172961 95069 172989
rect 95103 172961 95131 172989
rect 18117 164147 18145 164175
rect 18179 164147 18207 164175
rect 18241 164147 18269 164175
rect 18303 164147 18331 164175
rect 18117 164085 18145 164113
rect 18179 164085 18207 164113
rect 18241 164085 18269 164113
rect 18303 164085 18331 164113
rect 18117 164023 18145 164051
rect 18179 164023 18207 164051
rect 18241 164023 18269 164051
rect 18303 164023 18331 164051
rect 18117 163961 18145 163989
rect 18179 163961 18207 163989
rect 18241 163961 18269 163989
rect 18303 163961 18331 163989
rect 18117 155147 18145 155175
rect 18179 155147 18207 155175
rect 18241 155147 18269 155175
rect 18303 155147 18331 155175
rect 18117 155085 18145 155113
rect 18179 155085 18207 155113
rect 18241 155085 18269 155113
rect 18303 155085 18331 155113
rect 18117 155023 18145 155051
rect 18179 155023 18207 155051
rect 18241 155023 18269 155051
rect 18303 155023 18331 155051
rect 18117 154961 18145 154989
rect 18179 154961 18207 154989
rect 18241 154961 18269 154989
rect 18303 154961 18331 154989
rect 18117 146147 18145 146175
rect 18179 146147 18207 146175
rect 18241 146147 18269 146175
rect 18303 146147 18331 146175
rect 18117 146085 18145 146113
rect 18179 146085 18207 146113
rect 18241 146085 18269 146113
rect 18303 146085 18331 146113
rect 18117 146023 18145 146051
rect 18179 146023 18207 146051
rect 18241 146023 18269 146051
rect 18303 146023 18331 146051
rect 18117 145961 18145 145989
rect 18179 145961 18207 145989
rect 18241 145961 18269 145989
rect 18303 145961 18331 145989
rect 4617 140147 4645 140175
rect 4679 140147 4707 140175
rect 4741 140147 4769 140175
rect 4803 140147 4831 140175
rect 4617 140085 4645 140113
rect 4679 140085 4707 140113
rect 4741 140085 4769 140113
rect 4803 140085 4831 140113
rect 4617 140023 4645 140051
rect 4679 140023 4707 140051
rect 4741 140023 4769 140051
rect 4803 140023 4831 140051
rect 4617 139961 4645 139989
rect 4679 139961 4707 139989
rect 4741 139961 4769 139989
rect 4803 139961 4831 139989
rect 2757 38147 2785 38175
rect 2819 38147 2847 38175
rect 2881 38147 2909 38175
rect 2943 38147 2971 38175
rect 2757 38085 2785 38113
rect 2819 38085 2847 38113
rect 2881 38085 2909 38113
rect 2943 38085 2971 38113
rect 2757 38023 2785 38051
rect 2819 38023 2847 38051
rect 2881 38023 2909 38051
rect 2943 38023 2971 38051
rect 2757 37961 2785 37989
rect 2819 37961 2847 37989
rect 2881 37961 2909 37989
rect 2943 37961 2971 37989
rect 2757 29147 2785 29175
rect 2819 29147 2847 29175
rect 2881 29147 2909 29175
rect 2943 29147 2971 29175
rect 2757 29085 2785 29113
rect 2819 29085 2847 29113
rect 2881 29085 2909 29113
rect 2943 29085 2971 29113
rect 2757 29023 2785 29051
rect 2819 29023 2847 29051
rect 2881 29023 2909 29051
rect 2943 29023 2971 29051
rect 2757 28961 2785 28989
rect 2819 28961 2847 28989
rect 2881 28961 2909 28989
rect 2943 28961 2971 28989
rect 2757 20147 2785 20175
rect 2819 20147 2847 20175
rect 2881 20147 2909 20175
rect 2943 20147 2971 20175
rect 2757 20085 2785 20113
rect 2819 20085 2847 20113
rect 2881 20085 2909 20113
rect 2943 20085 2971 20113
rect 2757 20023 2785 20051
rect 2819 20023 2847 20051
rect 2881 20023 2909 20051
rect 2943 20023 2971 20051
rect 2757 19961 2785 19989
rect 2819 19961 2847 19989
rect 2881 19961 2909 19989
rect 2943 19961 2971 19989
rect 4617 131147 4645 131175
rect 4679 131147 4707 131175
rect 4741 131147 4769 131175
rect 4803 131147 4831 131175
rect 4617 131085 4645 131113
rect 4679 131085 4707 131113
rect 4741 131085 4769 131113
rect 4803 131085 4831 131113
rect 4617 131023 4645 131051
rect 4679 131023 4707 131051
rect 4741 131023 4769 131051
rect 4803 131023 4831 131051
rect 4617 130961 4645 130989
rect 4679 130961 4707 130989
rect 4741 130961 4769 130989
rect 4803 130961 4831 130989
rect 4617 122147 4645 122175
rect 4679 122147 4707 122175
rect 4741 122147 4769 122175
rect 4803 122147 4831 122175
rect 4617 122085 4645 122113
rect 4679 122085 4707 122113
rect 4741 122085 4769 122113
rect 4803 122085 4831 122113
rect 4617 122023 4645 122051
rect 4679 122023 4707 122051
rect 4741 122023 4769 122051
rect 4803 122023 4831 122051
rect 4617 121961 4645 121989
rect 4679 121961 4707 121989
rect 4741 121961 4769 121989
rect 4803 121961 4831 121989
rect 4617 113147 4645 113175
rect 4679 113147 4707 113175
rect 4741 113147 4769 113175
rect 4803 113147 4831 113175
rect 4617 113085 4645 113113
rect 4679 113085 4707 113113
rect 4741 113085 4769 113113
rect 4803 113085 4831 113113
rect 4617 113023 4645 113051
rect 4679 113023 4707 113051
rect 4741 113023 4769 113051
rect 4803 113023 4831 113051
rect 4617 112961 4645 112989
rect 4679 112961 4707 112989
rect 4741 112961 4769 112989
rect 4803 112961 4831 112989
rect 4617 104147 4645 104175
rect 4679 104147 4707 104175
rect 4741 104147 4769 104175
rect 4803 104147 4831 104175
rect 4617 104085 4645 104113
rect 4679 104085 4707 104113
rect 4741 104085 4769 104113
rect 4803 104085 4831 104113
rect 4617 104023 4645 104051
rect 4679 104023 4707 104051
rect 4741 104023 4769 104051
rect 4803 104023 4831 104051
rect 4617 103961 4645 103989
rect 4679 103961 4707 103989
rect 4741 103961 4769 103989
rect 4803 103961 4831 103989
rect 4617 95147 4645 95175
rect 4679 95147 4707 95175
rect 4741 95147 4769 95175
rect 4803 95147 4831 95175
rect 4617 95085 4645 95113
rect 4679 95085 4707 95113
rect 4741 95085 4769 95113
rect 4803 95085 4831 95113
rect 4617 95023 4645 95051
rect 4679 95023 4707 95051
rect 4741 95023 4769 95051
rect 4803 95023 4831 95051
rect 4617 94961 4645 94989
rect 4679 94961 4707 94989
rect 4741 94961 4769 94989
rect 4803 94961 4831 94989
rect 4617 86147 4645 86175
rect 4679 86147 4707 86175
rect 4741 86147 4769 86175
rect 4803 86147 4831 86175
rect 4617 86085 4645 86113
rect 4679 86085 4707 86113
rect 4741 86085 4769 86113
rect 4803 86085 4831 86113
rect 4617 86023 4645 86051
rect 4679 86023 4707 86051
rect 4741 86023 4769 86051
rect 4803 86023 4831 86051
rect 4617 85961 4645 85989
rect 4679 85961 4707 85989
rect 4741 85961 4769 85989
rect 4803 85961 4831 85989
rect 4617 77147 4645 77175
rect 4679 77147 4707 77175
rect 4741 77147 4769 77175
rect 4803 77147 4831 77175
rect 4617 77085 4645 77113
rect 4679 77085 4707 77113
rect 4741 77085 4769 77113
rect 4803 77085 4831 77113
rect 4617 77023 4645 77051
rect 4679 77023 4707 77051
rect 4741 77023 4769 77051
rect 4803 77023 4831 77051
rect 4617 76961 4645 76989
rect 4679 76961 4707 76989
rect 4741 76961 4769 76989
rect 4803 76961 4831 76989
rect 4617 68147 4645 68175
rect 4679 68147 4707 68175
rect 4741 68147 4769 68175
rect 4803 68147 4831 68175
rect 4617 68085 4645 68113
rect 4679 68085 4707 68113
rect 4741 68085 4769 68113
rect 4803 68085 4831 68113
rect 4617 68023 4645 68051
rect 4679 68023 4707 68051
rect 4741 68023 4769 68051
rect 4803 68023 4831 68051
rect 4617 67961 4645 67989
rect 4679 67961 4707 67989
rect 4741 67961 4769 67989
rect 4803 67961 4831 67989
rect 4617 59147 4645 59175
rect 4679 59147 4707 59175
rect 4741 59147 4769 59175
rect 4803 59147 4831 59175
rect 4617 59085 4645 59113
rect 4679 59085 4707 59113
rect 4741 59085 4769 59113
rect 4803 59085 4831 59113
rect 4617 59023 4645 59051
rect 4679 59023 4707 59051
rect 4741 59023 4769 59051
rect 4803 59023 4831 59051
rect 4617 58961 4645 58989
rect 4679 58961 4707 58989
rect 4741 58961 4769 58989
rect 4803 58961 4831 58989
rect 4617 50147 4645 50175
rect 4679 50147 4707 50175
rect 4741 50147 4769 50175
rect 4803 50147 4831 50175
rect 4617 50085 4645 50113
rect 4679 50085 4707 50113
rect 4741 50085 4769 50113
rect 4803 50085 4831 50113
rect 4617 50023 4645 50051
rect 4679 50023 4707 50051
rect 4741 50023 4769 50051
rect 4803 50023 4831 50051
rect 4617 49961 4645 49989
rect 4679 49961 4707 49989
rect 4741 49961 4769 49989
rect 4803 49961 4831 49989
rect 4617 41147 4645 41175
rect 4679 41147 4707 41175
rect 4741 41147 4769 41175
rect 4803 41147 4831 41175
rect 4617 41085 4645 41113
rect 4679 41085 4707 41113
rect 4741 41085 4769 41113
rect 4803 41085 4831 41113
rect 4617 41023 4645 41051
rect 4679 41023 4707 41051
rect 4741 41023 4769 41051
rect 4803 41023 4831 41051
rect 4617 40961 4645 40989
rect 4679 40961 4707 40989
rect 4741 40961 4769 40989
rect 4803 40961 4831 40989
rect 4617 32147 4645 32175
rect 4679 32147 4707 32175
rect 4741 32147 4769 32175
rect 4803 32147 4831 32175
rect 4617 32085 4645 32113
rect 4679 32085 4707 32113
rect 4741 32085 4769 32113
rect 4803 32085 4831 32113
rect 4617 32023 4645 32051
rect 4679 32023 4707 32051
rect 4741 32023 4769 32051
rect 4803 32023 4831 32051
rect 4617 31961 4645 31989
rect 4679 31961 4707 31989
rect 4741 31961 4769 31989
rect 4803 31961 4831 31989
rect 18117 137147 18145 137175
rect 18179 137147 18207 137175
rect 18241 137147 18269 137175
rect 18303 137147 18331 137175
rect 18117 137085 18145 137113
rect 18179 137085 18207 137113
rect 18241 137085 18269 137113
rect 18303 137085 18331 137113
rect 18117 137023 18145 137051
rect 18179 137023 18207 137051
rect 18241 137023 18269 137051
rect 18303 137023 18331 137051
rect 18117 136961 18145 136989
rect 18179 136961 18207 136989
rect 18241 136961 18269 136989
rect 18303 136961 18331 136989
rect 19977 167147 20005 167175
rect 20039 167147 20067 167175
rect 20101 167147 20129 167175
rect 20163 167147 20191 167175
rect 19977 167085 20005 167113
rect 20039 167085 20067 167113
rect 20101 167085 20129 167113
rect 20163 167085 20191 167113
rect 19977 167023 20005 167051
rect 20039 167023 20067 167051
rect 20101 167023 20129 167051
rect 20163 167023 20191 167051
rect 19977 166961 20005 166989
rect 20039 166961 20067 166989
rect 20101 166961 20129 166989
rect 20163 166961 20191 166989
rect 19977 158147 20005 158175
rect 20039 158147 20067 158175
rect 20101 158147 20129 158175
rect 20163 158147 20191 158175
rect 19977 158085 20005 158113
rect 20039 158085 20067 158113
rect 20101 158085 20129 158113
rect 20163 158085 20191 158113
rect 19977 158023 20005 158051
rect 20039 158023 20067 158051
rect 20101 158023 20129 158051
rect 20163 158023 20191 158051
rect 19977 157961 20005 157989
rect 20039 157961 20067 157989
rect 20101 157961 20129 157989
rect 20163 157961 20191 157989
rect 33477 164147 33505 164175
rect 33539 164147 33567 164175
rect 33601 164147 33629 164175
rect 33663 164147 33691 164175
rect 33477 164085 33505 164113
rect 33539 164085 33567 164113
rect 33601 164085 33629 164113
rect 33663 164085 33691 164113
rect 33477 164023 33505 164051
rect 33539 164023 33567 164051
rect 33601 164023 33629 164051
rect 33663 164023 33691 164051
rect 33477 163961 33505 163989
rect 33539 163961 33567 163989
rect 33601 163961 33629 163989
rect 33663 163961 33691 163989
rect 32259 155147 32287 155175
rect 32321 155147 32349 155175
rect 32259 155085 32287 155113
rect 32321 155085 32349 155113
rect 32259 155023 32287 155051
rect 32321 155023 32349 155051
rect 32259 154961 32287 154989
rect 32321 154961 32349 154989
rect 33477 155147 33505 155175
rect 33539 155147 33567 155175
rect 33601 155147 33629 155175
rect 33663 155147 33691 155175
rect 33477 155085 33505 155113
rect 33539 155085 33567 155113
rect 33601 155085 33629 155113
rect 33663 155085 33691 155113
rect 33477 155023 33505 155051
rect 33539 155023 33567 155051
rect 33601 155023 33629 155051
rect 33663 155023 33691 155051
rect 33477 154961 33505 154989
rect 33539 154961 33567 154989
rect 33601 154961 33629 154989
rect 33663 154961 33691 154989
rect 19977 149147 20005 149175
rect 20039 149147 20067 149175
rect 20101 149147 20129 149175
rect 20163 149147 20191 149175
rect 19977 149085 20005 149113
rect 20039 149085 20067 149113
rect 20101 149085 20129 149113
rect 20163 149085 20191 149113
rect 19977 149023 20005 149051
rect 20039 149023 20067 149051
rect 20101 149023 20129 149051
rect 20163 149023 20191 149051
rect 19977 148961 20005 148989
rect 20039 148961 20067 148989
rect 20101 148961 20129 148989
rect 20163 148961 20191 148989
rect 32259 146147 32287 146175
rect 32321 146147 32349 146175
rect 32259 146085 32287 146113
rect 32321 146085 32349 146113
rect 32259 146023 32287 146051
rect 32321 146023 32349 146051
rect 32259 145961 32287 145989
rect 32321 145961 32349 145989
rect 33477 146147 33505 146175
rect 33539 146147 33567 146175
rect 33601 146147 33629 146175
rect 33663 146147 33691 146175
rect 33477 146085 33505 146113
rect 33539 146085 33567 146113
rect 33601 146085 33629 146113
rect 33663 146085 33691 146113
rect 33477 146023 33505 146051
rect 33539 146023 33567 146051
rect 33601 146023 33629 146051
rect 33663 146023 33691 146051
rect 33477 145961 33505 145989
rect 33539 145961 33567 145989
rect 33601 145961 33629 145989
rect 33663 145961 33691 145989
rect 19977 140147 20005 140175
rect 20039 140147 20067 140175
rect 20101 140147 20129 140175
rect 20163 140147 20191 140175
rect 19977 140085 20005 140113
rect 20039 140085 20067 140113
rect 20101 140085 20129 140113
rect 20163 140085 20191 140113
rect 19977 140023 20005 140051
rect 20039 140023 20067 140051
rect 20101 140023 20129 140051
rect 20163 140023 20191 140051
rect 19977 139961 20005 139989
rect 20039 139961 20067 139989
rect 20101 139961 20129 139989
rect 20163 139961 20191 139989
rect 18117 128147 18145 128175
rect 18179 128147 18207 128175
rect 18241 128147 18269 128175
rect 18303 128147 18331 128175
rect 18117 128085 18145 128113
rect 18179 128085 18207 128113
rect 18241 128085 18269 128113
rect 18303 128085 18331 128113
rect 18117 128023 18145 128051
rect 18179 128023 18207 128051
rect 18241 128023 18269 128051
rect 18303 128023 18331 128051
rect 18117 127961 18145 127989
rect 18179 127961 18207 127989
rect 18241 127961 18269 127989
rect 18303 127961 18331 127989
rect 18117 119147 18145 119175
rect 18179 119147 18207 119175
rect 18241 119147 18269 119175
rect 18303 119147 18331 119175
rect 18117 119085 18145 119113
rect 18179 119085 18207 119113
rect 18241 119085 18269 119113
rect 18303 119085 18331 119113
rect 18117 119023 18145 119051
rect 18179 119023 18207 119051
rect 18241 119023 18269 119051
rect 18303 119023 18331 119051
rect 18117 118961 18145 118989
rect 18179 118961 18207 118989
rect 18241 118961 18269 118989
rect 18303 118961 18331 118989
rect 18117 110147 18145 110175
rect 18179 110147 18207 110175
rect 18241 110147 18269 110175
rect 18303 110147 18331 110175
rect 18117 110085 18145 110113
rect 18179 110085 18207 110113
rect 18241 110085 18269 110113
rect 18303 110085 18331 110113
rect 18117 110023 18145 110051
rect 18179 110023 18207 110051
rect 18241 110023 18269 110051
rect 18303 110023 18331 110051
rect 18117 109961 18145 109989
rect 18179 109961 18207 109989
rect 18241 109961 18269 109989
rect 18303 109961 18331 109989
rect 16259 101147 16287 101175
rect 16321 101147 16349 101175
rect 16259 101085 16287 101113
rect 16321 101085 16349 101113
rect 16259 101023 16287 101051
rect 16321 101023 16349 101051
rect 16259 100961 16287 100989
rect 16321 100961 16349 100989
rect 18117 101147 18145 101175
rect 18179 101147 18207 101175
rect 18241 101147 18269 101175
rect 18303 101147 18331 101175
rect 18117 101085 18145 101113
rect 18179 101085 18207 101113
rect 18241 101085 18269 101113
rect 18303 101085 18331 101113
rect 18117 101023 18145 101051
rect 18179 101023 18207 101051
rect 18241 101023 18269 101051
rect 18303 101023 18331 101051
rect 18117 100961 18145 100989
rect 18179 100961 18207 100989
rect 18241 100961 18269 100989
rect 18303 100961 18331 100989
rect 16259 92147 16287 92175
rect 16321 92147 16349 92175
rect 16259 92085 16287 92113
rect 16321 92085 16349 92113
rect 16259 92023 16287 92051
rect 16321 92023 16349 92051
rect 16259 91961 16287 91989
rect 16321 91961 16349 91989
rect 18117 92147 18145 92175
rect 18179 92147 18207 92175
rect 18241 92147 18269 92175
rect 18303 92147 18331 92175
rect 18117 92085 18145 92113
rect 18179 92085 18207 92113
rect 18241 92085 18269 92113
rect 18303 92085 18331 92113
rect 18117 92023 18145 92051
rect 18179 92023 18207 92051
rect 18241 92023 18269 92051
rect 18303 92023 18331 92051
rect 18117 91961 18145 91989
rect 18179 91961 18207 91989
rect 18241 91961 18269 91989
rect 18303 91961 18331 91989
rect 16259 83147 16287 83175
rect 16321 83147 16349 83175
rect 16259 83085 16287 83113
rect 16321 83085 16349 83113
rect 16259 83023 16287 83051
rect 16321 83023 16349 83051
rect 16259 82961 16287 82989
rect 16321 82961 16349 82989
rect 18117 83147 18145 83175
rect 18179 83147 18207 83175
rect 18241 83147 18269 83175
rect 18303 83147 18331 83175
rect 18117 83085 18145 83113
rect 18179 83085 18207 83113
rect 18241 83085 18269 83113
rect 18303 83085 18331 83113
rect 18117 83023 18145 83051
rect 18179 83023 18207 83051
rect 18241 83023 18269 83051
rect 18303 83023 18331 83051
rect 18117 82961 18145 82989
rect 18179 82961 18207 82989
rect 18241 82961 18269 82989
rect 18303 82961 18331 82989
rect 19977 131147 20005 131175
rect 20039 131147 20067 131175
rect 20101 131147 20129 131175
rect 20163 131147 20191 131175
rect 19977 131085 20005 131113
rect 20039 131085 20067 131113
rect 20101 131085 20129 131113
rect 20163 131085 20191 131113
rect 19977 131023 20005 131051
rect 20039 131023 20067 131051
rect 20101 131023 20129 131051
rect 20163 131023 20191 131051
rect 19977 130961 20005 130989
rect 20039 130961 20067 130989
rect 20101 130961 20129 130989
rect 20163 130961 20191 130989
rect 19977 122147 20005 122175
rect 20039 122147 20067 122175
rect 20101 122147 20129 122175
rect 20163 122147 20191 122175
rect 19977 122085 20005 122113
rect 20039 122085 20067 122113
rect 20101 122085 20129 122113
rect 20163 122085 20191 122113
rect 19977 122023 20005 122051
rect 20039 122023 20067 122051
rect 20101 122023 20129 122051
rect 20163 122023 20191 122051
rect 19977 121961 20005 121989
rect 20039 121961 20067 121989
rect 20101 121961 20129 121989
rect 20163 121961 20191 121989
rect 19977 113147 20005 113175
rect 20039 113147 20067 113175
rect 20101 113147 20129 113175
rect 20163 113147 20191 113175
rect 19977 113085 20005 113113
rect 20039 113085 20067 113113
rect 20101 113085 20129 113113
rect 20163 113085 20191 113113
rect 19977 113023 20005 113051
rect 20039 113023 20067 113051
rect 20101 113023 20129 113051
rect 20163 113023 20191 113051
rect 19977 112961 20005 112989
rect 20039 112961 20067 112989
rect 20101 112961 20129 112989
rect 20163 112961 20191 112989
rect 19977 104147 20005 104175
rect 20039 104147 20067 104175
rect 20101 104147 20129 104175
rect 20163 104147 20191 104175
rect 19977 104085 20005 104113
rect 20039 104085 20067 104113
rect 20101 104085 20129 104113
rect 20163 104085 20191 104113
rect 19977 104023 20005 104051
rect 20039 104023 20067 104051
rect 20101 104023 20129 104051
rect 20163 104023 20191 104051
rect 19977 103961 20005 103989
rect 20039 103961 20067 103989
rect 20101 103961 20129 103989
rect 20163 103961 20191 103989
rect 19977 95147 20005 95175
rect 20039 95147 20067 95175
rect 20101 95147 20129 95175
rect 20163 95147 20191 95175
rect 19977 95085 20005 95113
rect 20039 95085 20067 95113
rect 20101 95085 20129 95113
rect 20163 95085 20191 95113
rect 19977 95023 20005 95051
rect 20039 95023 20067 95051
rect 20101 95023 20129 95051
rect 20163 95023 20191 95051
rect 19977 94961 20005 94989
rect 20039 94961 20067 94989
rect 20101 94961 20129 94989
rect 20163 94961 20191 94989
rect 19977 86147 20005 86175
rect 20039 86147 20067 86175
rect 20101 86147 20129 86175
rect 20163 86147 20191 86175
rect 19977 86085 20005 86113
rect 20039 86085 20067 86113
rect 20101 86085 20129 86113
rect 20163 86085 20191 86113
rect 19977 86023 20005 86051
rect 20039 86023 20067 86051
rect 20101 86023 20129 86051
rect 20163 86023 20191 86051
rect 19977 85961 20005 85989
rect 20039 85961 20067 85989
rect 20101 85961 20129 85989
rect 20163 85961 20191 85989
rect 19977 77147 20005 77175
rect 20039 77147 20067 77175
rect 20101 77147 20129 77175
rect 20163 77147 20191 77175
rect 19977 77085 20005 77113
rect 20039 77085 20067 77113
rect 20101 77085 20129 77113
rect 20163 77085 20191 77113
rect 19977 77023 20005 77051
rect 20039 77023 20067 77051
rect 20101 77023 20129 77051
rect 20163 77023 20191 77051
rect 19977 76961 20005 76989
rect 20039 76961 20067 76989
rect 20101 76961 20129 76989
rect 20163 76961 20191 76989
rect 18117 74147 18145 74175
rect 18179 74147 18207 74175
rect 18241 74147 18269 74175
rect 18303 74147 18331 74175
rect 18117 74085 18145 74113
rect 18179 74085 18207 74113
rect 18241 74085 18269 74113
rect 18303 74085 18331 74113
rect 18117 74023 18145 74051
rect 18179 74023 18207 74051
rect 18241 74023 18269 74051
rect 18303 74023 18331 74051
rect 18117 73961 18145 73989
rect 18179 73961 18207 73989
rect 18241 73961 18269 73989
rect 18303 73961 18331 73989
rect 18117 65147 18145 65175
rect 18179 65147 18207 65175
rect 18241 65147 18269 65175
rect 18303 65147 18331 65175
rect 18117 65085 18145 65113
rect 18179 65085 18207 65113
rect 18241 65085 18269 65113
rect 18303 65085 18331 65113
rect 18117 65023 18145 65051
rect 18179 65023 18207 65051
rect 18241 65023 18269 65051
rect 18303 65023 18331 65051
rect 18117 64961 18145 64989
rect 18179 64961 18207 64989
rect 18241 64961 18269 64989
rect 18303 64961 18331 64989
rect 18117 56147 18145 56175
rect 18179 56147 18207 56175
rect 18241 56147 18269 56175
rect 18303 56147 18331 56175
rect 18117 56085 18145 56113
rect 18179 56085 18207 56113
rect 18241 56085 18269 56113
rect 18303 56085 18331 56113
rect 18117 56023 18145 56051
rect 18179 56023 18207 56051
rect 18241 56023 18269 56051
rect 18303 56023 18331 56051
rect 18117 55961 18145 55989
rect 18179 55961 18207 55989
rect 18241 55961 18269 55989
rect 18303 55961 18331 55989
rect 18117 47147 18145 47175
rect 18179 47147 18207 47175
rect 18241 47147 18269 47175
rect 18303 47147 18331 47175
rect 18117 47085 18145 47113
rect 18179 47085 18207 47113
rect 18241 47085 18269 47113
rect 18303 47085 18331 47113
rect 18117 47023 18145 47051
rect 18179 47023 18207 47051
rect 18241 47023 18269 47051
rect 18303 47023 18331 47051
rect 18117 46961 18145 46989
rect 18179 46961 18207 46989
rect 18241 46961 18269 46989
rect 18303 46961 18331 46989
rect 18117 38147 18145 38175
rect 18179 38147 18207 38175
rect 18241 38147 18269 38175
rect 18303 38147 18331 38175
rect 18117 38085 18145 38113
rect 18179 38085 18207 38113
rect 18241 38085 18269 38113
rect 18303 38085 18331 38113
rect 18117 38023 18145 38051
rect 18179 38023 18207 38051
rect 18241 38023 18269 38051
rect 18303 38023 18331 38051
rect 18117 37961 18145 37989
rect 18179 37961 18207 37989
rect 18241 37961 18269 37989
rect 18303 37961 18331 37989
rect 18117 29147 18145 29175
rect 18179 29147 18207 29175
rect 18241 29147 18269 29175
rect 18303 29147 18331 29175
rect 18117 29085 18145 29113
rect 18179 29085 18207 29113
rect 18241 29085 18269 29113
rect 18303 29085 18331 29113
rect 18117 29023 18145 29051
rect 18179 29023 18207 29051
rect 18241 29023 18269 29051
rect 18303 29023 18331 29051
rect 18117 28961 18145 28989
rect 18179 28961 18207 28989
rect 18241 28961 18269 28989
rect 18303 28961 18331 28989
rect 4617 23147 4645 23175
rect 4679 23147 4707 23175
rect 4741 23147 4769 23175
rect 4803 23147 4831 23175
rect 4617 23085 4645 23113
rect 4679 23085 4707 23113
rect 4741 23085 4769 23113
rect 4803 23085 4831 23113
rect 4617 23023 4645 23051
rect 4679 23023 4707 23051
rect 4741 23023 4769 23051
rect 4803 23023 4831 23051
rect 4617 22961 4645 22989
rect 4679 22961 4707 22989
rect 4741 22961 4769 22989
rect 4803 22961 4831 22989
rect 2757 11147 2785 11175
rect 2819 11147 2847 11175
rect 2881 11147 2909 11175
rect 2943 11147 2971 11175
rect 2757 11085 2785 11113
rect 2819 11085 2847 11113
rect 2881 11085 2909 11113
rect 2943 11085 2971 11113
rect 2757 11023 2785 11051
rect 2819 11023 2847 11051
rect 2881 11023 2909 11051
rect 2943 11023 2971 11051
rect 2757 10961 2785 10989
rect 2819 10961 2847 10989
rect 2881 10961 2909 10989
rect 2943 10961 2971 10989
rect -430 2147 -402 2175
rect -368 2147 -340 2175
rect -306 2147 -278 2175
rect -244 2147 -216 2175
rect -430 2085 -402 2113
rect -368 2085 -340 2113
rect -306 2085 -278 2113
rect -244 2085 -216 2113
rect -430 2023 -402 2051
rect -368 2023 -340 2051
rect -306 2023 -278 2051
rect -244 2023 -216 2051
rect -430 1961 -402 1989
rect -368 1961 -340 1989
rect -306 1961 -278 1989
rect -244 1961 -216 1989
rect -430 -108 -402 -80
rect -368 -108 -340 -80
rect -306 -108 -278 -80
rect -244 -108 -216 -80
rect -430 -170 -402 -142
rect -368 -170 -340 -142
rect -306 -170 -278 -142
rect -244 -170 -216 -142
rect -430 -232 -402 -204
rect -368 -232 -340 -204
rect -306 -232 -278 -204
rect -244 -232 -216 -204
rect -430 -294 -402 -266
rect -368 -294 -340 -266
rect -306 -294 -278 -266
rect -244 -294 -216 -266
rect 2757 2147 2785 2175
rect 2819 2147 2847 2175
rect 2881 2147 2909 2175
rect 2943 2147 2971 2175
rect 2757 2085 2785 2113
rect 2819 2085 2847 2113
rect 2881 2085 2909 2113
rect 2943 2085 2971 2113
rect 2757 2023 2785 2051
rect 2819 2023 2847 2051
rect 2881 2023 2909 2051
rect 2943 2023 2971 2051
rect 2757 1961 2785 1989
rect 2819 1961 2847 1989
rect 2881 1961 2909 1989
rect 2943 1961 2971 1989
rect 2757 -108 2785 -80
rect 2819 -108 2847 -80
rect 2881 -108 2909 -80
rect 2943 -108 2971 -80
rect 2757 -170 2785 -142
rect 2819 -170 2847 -142
rect 2881 -170 2909 -142
rect 2943 -170 2971 -142
rect 2757 -232 2785 -204
rect 2819 -232 2847 -204
rect 2881 -232 2909 -204
rect 2943 -232 2971 -204
rect 2757 -294 2785 -266
rect 2819 -294 2847 -266
rect 2881 -294 2909 -266
rect 2943 -294 2971 -266
rect -910 -588 -882 -560
rect -848 -588 -820 -560
rect -786 -588 -758 -560
rect -724 -588 -696 -560
rect -910 -650 -882 -622
rect -848 -650 -820 -622
rect -786 -650 -758 -622
rect -724 -650 -696 -622
rect -910 -712 -882 -684
rect -848 -712 -820 -684
rect -786 -712 -758 -684
rect -724 -712 -696 -684
rect -910 -774 -882 -746
rect -848 -774 -820 -746
rect -786 -774 -758 -746
rect -724 -774 -696 -746
rect 4617 14147 4645 14175
rect 4679 14147 4707 14175
rect 4741 14147 4769 14175
rect 4803 14147 4831 14175
rect 4617 14085 4645 14113
rect 4679 14085 4707 14113
rect 4741 14085 4769 14113
rect 4803 14085 4831 14113
rect 4617 14023 4645 14051
rect 4679 14023 4707 14051
rect 4741 14023 4769 14051
rect 4803 14023 4831 14051
rect 4617 13961 4645 13989
rect 4679 13961 4707 13989
rect 4741 13961 4769 13989
rect 4803 13961 4831 13989
rect 4617 5147 4645 5175
rect 4679 5147 4707 5175
rect 4741 5147 4769 5175
rect 4803 5147 4831 5175
rect 4617 5085 4645 5113
rect 4679 5085 4707 5113
rect 4741 5085 4769 5113
rect 4803 5085 4831 5113
rect 4617 5023 4645 5051
rect 4679 5023 4707 5051
rect 4741 5023 4769 5051
rect 4803 5023 4831 5051
rect 4617 4961 4645 4989
rect 4679 4961 4707 4989
rect 4741 4961 4769 4989
rect 4803 4961 4831 4989
rect 4617 -588 4645 -560
rect 4679 -588 4707 -560
rect 4741 -588 4769 -560
rect 4803 -588 4831 -560
rect 4617 -650 4645 -622
rect 4679 -650 4707 -622
rect 4741 -650 4769 -622
rect 4803 -650 4831 -622
rect 4617 -712 4645 -684
rect 4679 -712 4707 -684
rect 4741 -712 4769 -684
rect 4803 -712 4831 -684
rect 4617 -774 4645 -746
rect 4679 -774 4707 -746
rect 4741 -774 4769 -746
rect 4803 -774 4831 -746
rect 18117 20147 18145 20175
rect 18179 20147 18207 20175
rect 18241 20147 18269 20175
rect 18303 20147 18331 20175
rect 18117 20085 18145 20113
rect 18179 20085 18207 20113
rect 18241 20085 18269 20113
rect 18303 20085 18331 20113
rect 18117 20023 18145 20051
rect 18179 20023 18207 20051
rect 18241 20023 18269 20051
rect 18303 20023 18331 20051
rect 18117 19961 18145 19989
rect 18179 19961 18207 19989
rect 18241 19961 18269 19989
rect 18303 19961 18331 19989
rect 18117 11147 18145 11175
rect 18179 11147 18207 11175
rect 18241 11147 18269 11175
rect 18303 11147 18331 11175
rect 18117 11085 18145 11113
rect 18179 11085 18207 11113
rect 18241 11085 18269 11113
rect 18303 11085 18331 11113
rect 18117 11023 18145 11051
rect 18179 11023 18207 11051
rect 18241 11023 18269 11051
rect 18303 11023 18331 11051
rect 18117 10961 18145 10989
rect 18179 10961 18207 10989
rect 18241 10961 18269 10989
rect 18303 10961 18331 10989
rect 18117 2147 18145 2175
rect 18179 2147 18207 2175
rect 18241 2147 18269 2175
rect 18303 2147 18331 2175
rect 18117 2085 18145 2113
rect 18179 2085 18207 2113
rect 18241 2085 18269 2113
rect 18303 2085 18331 2113
rect 18117 2023 18145 2051
rect 18179 2023 18207 2051
rect 18241 2023 18269 2051
rect 18303 2023 18331 2051
rect 18117 1961 18145 1989
rect 18179 1961 18207 1989
rect 18241 1961 18269 1989
rect 18303 1961 18331 1989
rect 18117 -108 18145 -80
rect 18179 -108 18207 -80
rect 18241 -108 18269 -80
rect 18303 -108 18331 -80
rect 18117 -170 18145 -142
rect 18179 -170 18207 -142
rect 18241 -170 18269 -142
rect 18303 -170 18331 -142
rect 18117 -232 18145 -204
rect 18179 -232 18207 -204
rect 18241 -232 18269 -204
rect 18303 -232 18331 -204
rect 18117 -294 18145 -266
rect 18179 -294 18207 -266
rect 18241 -294 18269 -266
rect 18303 -294 18331 -266
rect 32259 137147 32287 137175
rect 32321 137147 32349 137175
rect 32259 137085 32287 137113
rect 32321 137085 32349 137113
rect 32259 137023 32287 137051
rect 32321 137023 32349 137051
rect 32259 136961 32287 136989
rect 32321 136961 32349 136989
rect 33477 137147 33505 137175
rect 33539 137147 33567 137175
rect 33601 137147 33629 137175
rect 33663 137147 33691 137175
rect 33477 137085 33505 137113
rect 33539 137085 33567 137113
rect 33601 137085 33629 137113
rect 33663 137085 33691 137113
rect 33477 137023 33505 137051
rect 33539 137023 33567 137051
rect 33601 137023 33629 137051
rect 33663 137023 33691 137051
rect 33477 136961 33505 136989
rect 33539 136961 33567 136989
rect 33601 136961 33629 136989
rect 33663 136961 33691 136989
rect 33477 128147 33505 128175
rect 33539 128147 33567 128175
rect 33601 128147 33629 128175
rect 33663 128147 33691 128175
rect 33477 128085 33505 128113
rect 33539 128085 33567 128113
rect 33601 128085 33629 128113
rect 33663 128085 33691 128113
rect 33477 128023 33505 128051
rect 33539 128023 33567 128051
rect 33601 128023 33629 128051
rect 33663 128023 33691 128051
rect 33477 127961 33505 127989
rect 33539 127961 33567 127989
rect 33601 127961 33629 127989
rect 33663 127961 33691 127989
rect 33477 119147 33505 119175
rect 33539 119147 33567 119175
rect 33601 119147 33629 119175
rect 33663 119147 33691 119175
rect 33477 119085 33505 119113
rect 33539 119085 33567 119113
rect 33601 119085 33629 119113
rect 33663 119085 33691 119113
rect 33477 119023 33505 119051
rect 33539 119023 33567 119051
rect 33601 119023 33629 119051
rect 33663 119023 33691 119051
rect 33477 118961 33505 118989
rect 33539 118961 33567 118989
rect 33601 118961 33629 118989
rect 33663 118961 33691 118989
rect 33477 110147 33505 110175
rect 33539 110147 33567 110175
rect 33601 110147 33629 110175
rect 33663 110147 33691 110175
rect 33477 110085 33505 110113
rect 33539 110085 33567 110113
rect 33601 110085 33629 110113
rect 33663 110085 33691 110113
rect 33477 110023 33505 110051
rect 33539 110023 33567 110051
rect 33601 110023 33629 110051
rect 33663 110023 33691 110051
rect 33477 109961 33505 109989
rect 33539 109961 33567 109989
rect 33601 109961 33629 109989
rect 33663 109961 33691 109989
rect 31619 101147 31647 101175
rect 31681 101147 31709 101175
rect 31619 101085 31647 101113
rect 31681 101085 31709 101113
rect 31619 101023 31647 101051
rect 31681 101023 31709 101051
rect 31619 100961 31647 100989
rect 31681 100961 31709 100989
rect 33477 101147 33505 101175
rect 33539 101147 33567 101175
rect 33601 101147 33629 101175
rect 33663 101147 33691 101175
rect 33477 101085 33505 101113
rect 33539 101085 33567 101113
rect 33601 101085 33629 101113
rect 33663 101085 33691 101113
rect 33477 101023 33505 101051
rect 33539 101023 33567 101051
rect 33601 101023 33629 101051
rect 33663 101023 33691 101051
rect 33477 100961 33505 100989
rect 33539 100961 33567 100989
rect 33601 100961 33629 100989
rect 33663 100961 33691 100989
rect 23939 95147 23967 95175
rect 24001 95147 24029 95175
rect 23939 95085 23967 95113
rect 24001 95085 24029 95113
rect 23939 95023 23967 95051
rect 24001 95023 24029 95051
rect 23939 94961 23967 94989
rect 24001 94961 24029 94989
rect 31619 92147 31647 92175
rect 31681 92147 31709 92175
rect 31619 92085 31647 92113
rect 31681 92085 31709 92113
rect 31619 92023 31647 92051
rect 31681 92023 31709 92051
rect 31619 91961 31647 91989
rect 31681 91961 31709 91989
rect 33477 92147 33505 92175
rect 33539 92147 33567 92175
rect 33601 92147 33629 92175
rect 33663 92147 33691 92175
rect 33477 92085 33505 92113
rect 33539 92085 33567 92113
rect 33601 92085 33629 92113
rect 33663 92085 33691 92113
rect 33477 92023 33505 92051
rect 33539 92023 33567 92051
rect 33601 92023 33629 92051
rect 33663 92023 33691 92051
rect 33477 91961 33505 91989
rect 33539 91961 33567 91989
rect 33601 91961 33629 91989
rect 33663 91961 33691 91989
rect 35337 167147 35365 167175
rect 35399 167147 35427 167175
rect 35461 167147 35489 167175
rect 35523 167147 35551 167175
rect 35337 167085 35365 167113
rect 35399 167085 35427 167113
rect 35461 167085 35489 167113
rect 35523 167085 35551 167113
rect 35337 167023 35365 167051
rect 35399 167023 35427 167051
rect 35461 167023 35489 167051
rect 35523 167023 35551 167051
rect 35337 166961 35365 166989
rect 35399 166961 35427 166989
rect 35461 166961 35489 166989
rect 35523 166961 35551 166989
rect 48837 164147 48865 164175
rect 48899 164147 48927 164175
rect 48961 164147 48989 164175
rect 49023 164147 49051 164175
rect 48837 164085 48865 164113
rect 48899 164085 48927 164113
rect 48961 164085 48989 164113
rect 49023 164085 49051 164113
rect 48837 164023 48865 164051
rect 48899 164023 48927 164051
rect 48961 164023 48989 164051
rect 49023 164023 49051 164051
rect 48837 163961 48865 163989
rect 48899 163961 48927 163989
rect 48961 163961 48989 163989
rect 49023 163961 49051 163989
rect 35337 158147 35365 158175
rect 35399 158147 35427 158175
rect 35461 158147 35489 158175
rect 35523 158147 35551 158175
rect 35337 158085 35365 158113
rect 35399 158085 35427 158113
rect 35461 158085 35489 158113
rect 35523 158085 35551 158113
rect 35337 158023 35365 158051
rect 35399 158023 35427 158051
rect 35461 158023 35489 158051
rect 35523 158023 35551 158051
rect 35337 157961 35365 157989
rect 35399 157961 35427 157989
rect 35461 157961 35489 157989
rect 35523 157961 35551 157989
rect 39939 158147 39967 158175
rect 40001 158147 40029 158175
rect 39939 158085 39967 158113
rect 40001 158085 40029 158113
rect 39939 158023 39967 158051
rect 40001 158023 40029 158051
rect 39939 157961 39967 157989
rect 40001 157961 40029 157989
rect 47619 155147 47647 155175
rect 47681 155147 47709 155175
rect 47619 155085 47647 155113
rect 47681 155085 47709 155113
rect 47619 155023 47647 155051
rect 47681 155023 47709 155051
rect 47619 154961 47647 154989
rect 47681 154961 47709 154989
rect 48837 155147 48865 155175
rect 48899 155147 48927 155175
rect 48961 155147 48989 155175
rect 49023 155147 49051 155175
rect 48837 155085 48865 155113
rect 48899 155085 48927 155113
rect 48961 155085 48989 155113
rect 49023 155085 49051 155113
rect 48837 155023 48865 155051
rect 48899 155023 48927 155051
rect 48961 155023 48989 155051
rect 49023 155023 49051 155051
rect 48837 154961 48865 154989
rect 48899 154961 48927 154989
rect 48961 154961 48989 154989
rect 49023 154961 49051 154989
rect 35337 149147 35365 149175
rect 35399 149147 35427 149175
rect 35461 149147 35489 149175
rect 35523 149147 35551 149175
rect 35337 149085 35365 149113
rect 35399 149085 35427 149113
rect 35461 149085 35489 149113
rect 35523 149085 35551 149113
rect 35337 149023 35365 149051
rect 35399 149023 35427 149051
rect 35461 149023 35489 149051
rect 35523 149023 35551 149051
rect 35337 148961 35365 148989
rect 35399 148961 35427 148989
rect 35461 148961 35489 148989
rect 35523 148961 35551 148989
rect 39939 149147 39967 149175
rect 40001 149147 40029 149175
rect 39939 149085 39967 149113
rect 40001 149085 40029 149113
rect 39939 149023 39967 149051
rect 40001 149023 40029 149051
rect 39939 148961 39967 148989
rect 40001 148961 40029 148989
rect 47619 146147 47647 146175
rect 47681 146147 47709 146175
rect 47619 146085 47647 146113
rect 47681 146085 47709 146113
rect 47619 146023 47647 146051
rect 47681 146023 47709 146051
rect 47619 145961 47647 145989
rect 47681 145961 47709 145989
rect 48837 146147 48865 146175
rect 48899 146147 48927 146175
rect 48961 146147 48989 146175
rect 49023 146147 49051 146175
rect 48837 146085 48865 146113
rect 48899 146085 48927 146113
rect 48961 146085 48989 146113
rect 49023 146085 49051 146113
rect 48837 146023 48865 146051
rect 48899 146023 48927 146051
rect 48961 146023 48989 146051
rect 49023 146023 49051 146051
rect 48837 145961 48865 145989
rect 48899 145961 48927 145989
rect 48961 145961 48989 145989
rect 49023 145961 49051 145989
rect 35337 140147 35365 140175
rect 35399 140147 35427 140175
rect 35461 140147 35489 140175
rect 35523 140147 35551 140175
rect 35337 140085 35365 140113
rect 35399 140085 35427 140113
rect 35461 140085 35489 140113
rect 35523 140085 35551 140113
rect 35337 140023 35365 140051
rect 35399 140023 35427 140051
rect 35461 140023 35489 140051
rect 35523 140023 35551 140051
rect 35337 139961 35365 139989
rect 35399 139961 35427 139989
rect 35461 139961 35489 139989
rect 35523 139961 35551 139989
rect 39939 140147 39967 140175
rect 40001 140147 40029 140175
rect 39939 140085 39967 140113
rect 40001 140085 40029 140113
rect 39939 140023 39967 140051
rect 40001 140023 40029 140051
rect 39939 139961 39967 139989
rect 40001 139961 40029 139989
rect 47619 137147 47647 137175
rect 47681 137147 47709 137175
rect 47619 137085 47647 137113
rect 47681 137085 47709 137113
rect 47619 137023 47647 137051
rect 47681 137023 47709 137051
rect 47619 136961 47647 136989
rect 47681 136961 47709 136989
rect 48837 137147 48865 137175
rect 48899 137147 48927 137175
rect 48961 137147 48989 137175
rect 49023 137147 49051 137175
rect 48837 137085 48865 137113
rect 48899 137085 48927 137113
rect 48961 137085 48989 137113
rect 49023 137085 49051 137113
rect 48837 137023 48865 137051
rect 48899 137023 48927 137051
rect 48961 137023 48989 137051
rect 49023 137023 49051 137051
rect 48837 136961 48865 136989
rect 48899 136961 48927 136989
rect 48961 136961 48989 136989
rect 49023 136961 49051 136989
rect 35337 131147 35365 131175
rect 35399 131147 35427 131175
rect 35461 131147 35489 131175
rect 35523 131147 35551 131175
rect 35337 131085 35365 131113
rect 35399 131085 35427 131113
rect 35461 131085 35489 131113
rect 35523 131085 35551 131113
rect 35337 131023 35365 131051
rect 35399 131023 35427 131051
rect 35461 131023 35489 131051
rect 35523 131023 35551 131051
rect 35337 130961 35365 130989
rect 35399 130961 35427 130989
rect 35461 130961 35489 130989
rect 35523 130961 35551 130989
rect 35337 122147 35365 122175
rect 35399 122147 35427 122175
rect 35461 122147 35489 122175
rect 35523 122147 35551 122175
rect 35337 122085 35365 122113
rect 35399 122085 35427 122113
rect 35461 122085 35489 122113
rect 35523 122085 35551 122113
rect 35337 122023 35365 122051
rect 35399 122023 35427 122051
rect 35461 122023 35489 122051
rect 35523 122023 35551 122051
rect 35337 121961 35365 121989
rect 35399 121961 35427 121989
rect 35461 121961 35489 121989
rect 35523 121961 35551 121989
rect 35337 113147 35365 113175
rect 35399 113147 35427 113175
rect 35461 113147 35489 113175
rect 35523 113147 35551 113175
rect 35337 113085 35365 113113
rect 35399 113085 35427 113113
rect 35461 113085 35489 113113
rect 35523 113085 35551 113113
rect 35337 113023 35365 113051
rect 35399 113023 35427 113051
rect 35461 113023 35489 113051
rect 35523 113023 35551 113051
rect 35337 112961 35365 112989
rect 35399 112961 35427 112989
rect 35461 112961 35489 112989
rect 35523 112961 35551 112989
rect 35337 104147 35365 104175
rect 35399 104147 35427 104175
rect 35461 104147 35489 104175
rect 35523 104147 35551 104175
rect 35337 104085 35365 104113
rect 35399 104085 35427 104113
rect 35461 104085 35489 104113
rect 35523 104085 35551 104113
rect 35337 104023 35365 104051
rect 35399 104023 35427 104051
rect 35461 104023 35489 104051
rect 35523 104023 35551 104051
rect 35337 103961 35365 103989
rect 35399 103961 35427 103989
rect 35461 103961 35489 103989
rect 35523 103961 35551 103989
rect 48837 128147 48865 128175
rect 48899 128147 48927 128175
rect 48961 128147 48989 128175
rect 49023 128147 49051 128175
rect 48837 128085 48865 128113
rect 48899 128085 48927 128113
rect 48961 128085 48989 128113
rect 49023 128085 49051 128113
rect 48837 128023 48865 128051
rect 48899 128023 48927 128051
rect 48961 128023 48989 128051
rect 49023 128023 49051 128051
rect 48837 127961 48865 127989
rect 48899 127961 48927 127989
rect 48961 127961 48989 127989
rect 49023 127961 49051 127989
rect 48837 119147 48865 119175
rect 48899 119147 48927 119175
rect 48961 119147 48989 119175
rect 49023 119147 49051 119175
rect 48837 119085 48865 119113
rect 48899 119085 48927 119113
rect 48961 119085 48989 119113
rect 49023 119085 49051 119113
rect 48837 119023 48865 119051
rect 48899 119023 48927 119051
rect 48961 119023 48989 119051
rect 49023 119023 49051 119051
rect 48837 118961 48865 118989
rect 48899 118961 48927 118989
rect 48961 118961 48989 118989
rect 49023 118961 49051 118989
rect 48837 110147 48865 110175
rect 48899 110147 48927 110175
rect 48961 110147 48989 110175
rect 49023 110147 49051 110175
rect 48837 110085 48865 110113
rect 48899 110085 48927 110113
rect 48961 110085 48989 110113
rect 49023 110085 49051 110113
rect 48837 110023 48865 110051
rect 48899 110023 48927 110051
rect 48961 110023 48989 110051
rect 49023 110023 49051 110051
rect 48837 109961 48865 109989
rect 48899 109961 48927 109989
rect 48961 109961 48989 109989
rect 49023 109961 49051 109989
rect 46979 101147 47007 101175
rect 47041 101147 47069 101175
rect 46979 101085 47007 101113
rect 47041 101085 47069 101113
rect 46979 101023 47007 101051
rect 47041 101023 47069 101051
rect 46979 100961 47007 100989
rect 47041 100961 47069 100989
rect 48837 101147 48865 101175
rect 48899 101147 48927 101175
rect 48961 101147 48989 101175
rect 49023 101147 49051 101175
rect 48837 101085 48865 101113
rect 48899 101085 48927 101113
rect 48961 101085 48989 101113
rect 49023 101085 49051 101113
rect 48837 101023 48865 101051
rect 48899 101023 48927 101051
rect 48961 101023 48989 101051
rect 49023 101023 49051 101051
rect 48837 100961 48865 100989
rect 48899 100961 48927 100989
rect 48961 100961 48989 100989
rect 49023 100961 49051 100989
rect 35337 95147 35365 95175
rect 35399 95147 35427 95175
rect 35461 95147 35489 95175
rect 35523 95147 35551 95175
rect 35337 95085 35365 95113
rect 35399 95085 35427 95113
rect 35461 95085 35489 95113
rect 35523 95085 35551 95113
rect 35337 95023 35365 95051
rect 35399 95023 35427 95051
rect 35461 95023 35489 95051
rect 35523 95023 35551 95051
rect 35337 94961 35365 94989
rect 35399 94961 35427 94989
rect 35461 94961 35489 94989
rect 35523 94961 35551 94989
rect 39299 95147 39327 95175
rect 39361 95147 39389 95175
rect 39299 95085 39327 95113
rect 39361 95085 39389 95113
rect 39299 95023 39327 95051
rect 39361 95023 39389 95051
rect 39299 94961 39327 94989
rect 39361 94961 39389 94989
rect 46979 92147 47007 92175
rect 47041 92147 47069 92175
rect 46979 92085 47007 92113
rect 47041 92085 47069 92113
rect 46979 92023 47007 92051
rect 47041 92023 47069 92051
rect 46979 91961 47007 91989
rect 47041 91961 47069 91989
rect 48837 92147 48865 92175
rect 48899 92147 48927 92175
rect 48961 92147 48989 92175
rect 49023 92147 49051 92175
rect 48837 92085 48865 92113
rect 48899 92085 48927 92113
rect 48961 92085 48989 92113
rect 49023 92085 49051 92113
rect 48837 92023 48865 92051
rect 48899 92023 48927 92051
rect 48961 92023 48989 92051
rect 49023 92023 49051 92051
rect 48837 91961 48865 91989
rect 48899 91961 48927 91989
rect 48961 91961 48989 91989
rect 49023 91961 49051 91989
rect 50697 167147 50725 167175
rect 50759 167147 50787 167175
rect 50821 167147 50849 167175
rect 50883 167147 50911 167175
rect 50697 167085 50725 167113
rect 50759 167085 50787 167113
rect 50821 167085 50849 167113
rect 50883 167085 50911 167113
rect 50697 167023 50725 167051
rect 50759 167023 50787 167051
rect 50821 167023 50849 167051
rect 50883 167023 50911 167051
rect 50697 166961 50725 166989
rect 50759 166961 50787 166989
rect 50821 166961 50849 166989
rect 50883 166961 50911 166989
rect 64197 164147 64225 164175
rect 64259 164147 64287 164175
rect 64321 164147 64349 164175
rect 64383 164147 64411 164175
rect 64197 164085 64225 164113
rect 64259 164085 64287 164113
rect 64321 164085 64349 164113
rect 64383 164085 64411 164113
rect 64197 164023 64225 164051
rect 64259 164023 64287 164051
rect 64321 164023 64349 164051
rect 64383 164023 64411 164051
rect 64197 163961 64225 163989
rect 64259 163961 64287 163989
rect 64321 163961 64349 163989
rect 64383 163961 64411 163989
rect 50697 158147 50725 158175
rect 50759 158147 50787 158175
rect 50821 158147 50849 158175
rect 50883 158147 50911 158175
rect 50697 158085 50725 158113
rect 50759 158085 50787 158113
rect 50821 158085 50849 158113
rect 50883 158085 50911 158113
rect 50697 158023 50725 158051
rect 50759 158023 50787 158051
rect 50821 158023 50849 158051
rect 50883 158023 50911 158051
rect 50697 157961 50725 157989
rect 50759 157961 50787 157989
rect 50821 157961 50849 157989
rect 50883 157961 50911 157989
rect 55299 158147 55327 158175
rect 55361 158147 55389 158175
rect 55299 158085 55327 158113
rect 55361 158085 55389 158113
rect 55299 158023 55327 158051
rect 55361 158023 55389 158051
rect 55299 157961 55327 157989
rect 55361 157961 55389 157989
rect 62979 155147 63007 155175
rect 63041 155147 63069 155175
rect 62979 155085 63007 155113
rect 63041 155085 63069 155113
rect 62979 155023 63007 155051
rect 63041 155023 63069 155051
rect 62979 154961 63007 154989
rect 63041 154961 63069 154989
rect 64197 155147 64225 155175
rect 64259 155147 64287 155175
rect 64321 155147 64349 155175
rect 64383 155147 64411 155175
rect 64197 155085 64225 155113
rect 64259 155085 64287 155113
rect 64321 155085 64349 155113
rect 64383 155085 64411 155113
rect 64197 155023 64225 155051
rect 64259 155023 64287 155051
rect 64321 155023 64349 155051
rect 64383 155023 64411 155051
rect 64197 154961 64225 154989
rect 64259 154961 64287 154989
rect 64321 154961 64349 154989
rect 64383 154961 64411 154989
rect 50697 149147 50725 149175
rect 50759 149147 50787 149175
rect 50821 149147 50849 149175
rect 50883 149147 50911 149175
rect 50697 149085 50725 149113
rect 50759 149085 50787 149113
rect 50821 149085 50849 149113
rect 50883 149085 50911 149113
rect 50697 149023 50725 149051
rect 50759 149023 50787 149051
rect 50821 149023 50849 149051
rect 50883 149023 50911 149051
rect 50697 148961 50725 148989
rect 50759 148961 50787 148989
rect 50821 148961 50849 148989
rect 50883 148961 50911 148989
rect 55299 149147 55327 149175
rect 55361 149147 55389 149175
rect 55299 149085 55327 149113
rect 55361 149085 55389 149113
rect 55299 149023 55327 149051
rect 55361 149023 55389 149051
rect 55299 148961 55327 148989
rect 55361 148961 55389 148989
rect 62979 146147 63007 146175
rect 63041 146147 63069 146175
rect 62979 146085 63007 146113
rect 63041 146085 63069 146113
rect 62979 146023 63007 146051
rect 63041 146023 63069 146051
rect 62979 145961 63007 145989
rect 63041 145961 63069 145989
rect 64197 146147 64225 146175
rect 64259 146147 64287 146175
rect 64321 146147 64349 146175
rect 64383 146147 64411 146175
rect 64197 146085 64225 146113
rect 64259 146085 64287 146113
rect 64321 146085 64349 146113
rect 64383 146085 64411 146113
rect 64197 146023 64225 146051
rect 64259 146023 64287 146051
rect 64321 146023 64349 146051
rect 64383 146023 64411 146051
rect 64197 145961 64225 145989
rect 64259 145961 64287 145989
rect 64321 145961 64349 145989
rect 64383 145961 64411 145989
rect 50697 140147 50725 140175
rect 50759 140147 50787 140175
rect 50821 140147 50849 140175
rect 50883 140147 50911 140175
rect 50697 140085 50725 140113
rect 50759 140085 50787 140113
rect 50821 140085 50849 140113
rect 50883 140085 50911 140113
rect 50697 140023 50725 140051
rect 50759 140023 50787 140051
rect 50821 140023 50849 140051
rect 50883 140023 50911 140051
rect 50697 139961 50725 139989
rect 50759 139961 50787 139989
rect 50821 139961 50849 139989
rect 50883 139961 50911 139989
rect 55299 140147 55327 140175
rect 55361 140147 55389 140175
rect 55299 140085 55327 140113
rect 55361 140085 55389 140113
rect 55299 140023 55327 140051
rect 55361 140023 55389 140051
rect 55299 139961 55327 139989
rect 55361 139961 55389 139989
rect 62979 137147 63007 137175
rect 63041 137147 63069 137175
rect 62979 137085 63007 137113
rect 63041 137085 63069 137113
rect 62979 137023 63007 137051
rect 63041 137023 63069 137051
rect 62979 136961 63007 136989
rect 63041 136961 63069 136989
rect 64197 137147 64225 137175
rect 64259 137147 64287 137175
rect 64321 137147 64349 137175
rect 64383 137147 64411 137175
rect 64197 137085 64225 137113
rect 64259 137085 64287 137113
rect 64321 137085 64349 137113
rect 64383 137085 64411 137113
rect 64197 137023 64225 137051
rect 64259 137023 64287 137051
rect 64321 137023 64349 137051
rect 64383 137023 64411 137051
rect 64197 136961 64225 136989
rect 64259 136961 64287 136989
rect 64321 136961 64349 136989
rect 64383 136961 64411 136989
rect 50697 131147 50725 131175
rect 50759 131147 50787 131175
rect 50821 131147 50849 131175
rect 50883 131147 50911 131175
rect 50697 131085 50725 131113
rect 50759 131085 50787 131113
rect 50821 131085 50849 131113
rect 50883 131085 50911 131113
rect 50697 131023 50725 131051
rect 50759 131023 50787 131051
rect 50821 131023 50849 131051
rect 50883 131023 50911 131051
rect 50697 130961 50725 130989
rect 50759 130961 50787 130989
rect 50821 130961 50849 130989
rect 50883 130961 50911 130989
rect 50697 122147 50725 122175
rect 50759 122147 50787 122175
rect 50821 122147 50849 122175
rect 50883 122147 50911 122175
rect 50697 122085 50725 122113
rect 50759 122085 50787 122113
rect 50821 122085 50849 122113
rect 50883 122085 50911 122113
rect 50697 122023 50725 122051
rect 50759 122023 50787 122051
rect 50821 122023 50849 122051
rect 50883 122023 50911 122051
rect 50697 121961 50725 121989
rect 50759 121961 50787 121989
rect 50821 121961 50849 121989
rect 50883 121961 50911 121989
rect 50697 113147 50725 113175
rect 50759 113147 50787 113175
rect 50821 113147 50849 113175
rect 50883 113147 50911 113175
rect 50697 113085 50725 113113
rect 50759 113085 50787 113113
rect 50821 113085 50849 113113
rect 50883 113085 50911 113113
rect 50697 113023 50725 113051
rect 50759 113023 50787 113051
rect 50821 113023 50849 113051
rect 50883 113023 50911 113051
rect 50697 112961 50725 112989
rect 50759 112961 50787 112989
rect 50821 112961 50849 112989
rect 50883 112961 50911 112989
rect 50697 104147 50725 104175
rect 50759 104147 50787 104175
rect 50821 104147 50849 104175
rect 50883 104147 50911 104175
rect 50697 104085 50725 104113
rect 50759 104085 50787 104113
rect 50821 104085 50849 104113
rect 50883 104085 50911 104113
rect 50697 104023 50725 104051
rect 50759 104023 50787 104051
rect 50821 104023 50849 104051
rect 50883 104023 50911 104051
rect 50697 103961 50725 103989
rect 50759 103961 50787 103989
rect 50821 103961 50849 103989
rect 50883 103961 50911 103989
rect 64197 128147 64225 128175
rect 64259 128147 64287 128175
rect 64321 128147 64349 128175
rect 64383 128147 64411 128175
rect 64197 128085 64225 128113
rect 64259 128085 64287 128113
rect 64321 128085 64349 128113
rect 64383 128085 64411 128113
rect 64197 128023 64225 128051
rect 64259 128023 64287 128051
rect 64321 128023 64349 128051
rect 64383 128023 64411 128051
rect 64197 127961 64225 127989
rect 64259 127961 64287 127989
rect 64321 127961 64349 127989
rect 64383 127961 64411 127989
rect 64197 119147 64225 119175
rect 64259 119147 64287 119175
rect 64321 119147 64349 119175
rect 64383 119147 64411 119175
rect 64197 119085 64225 119113
rect 64259 119085 64287 119113
rect 64321 119085 64349 119113
rect 64383 119085 64411 119113
rect 64197 119023 64225 119051
rect 64259 119023 64287 119051
rect 64321 119023 64349 119051
rect 64383 119023 64411 119051
rect 64197 118961 64225 118989
rect 64259 118961 64287 118989
rect 64321 118961 64349 118989
rect 64383 118961 64411 118989
rect 64197 110147 64225 110175
rect 64259 110147 64287 110175
rect 64321 110147 64349 110175
rect 64383 110147 64411 110175
rect 64197 110085 64225 110113
rect 64259 110085 64287 110113
rect 64321 110085 64349 110113
rect 64383 110085 64411 110113
rect 64197 110023 64225 110051
rect 64259 110023 64287 110051
rect 64321 110023 64349 110051
rect 64383 110023 64411 110051
rect 64197 109961 64225 109989
rect 64259 109961 64287 109989
rect 64321 109961 64349 109989
rect 64383 109961 64411 109989
rect 62339 101147 62367 101175
rect 62401 101147 62429 101175
rect 62339 101085 62367 101113
rect 62401 101085 62429 101113
rect 62339 101023 62367 101051
rect 62401 101023 62429 101051
rect 62339 100961 62367 100989
rect 62401 100961 62429 100989
rect 64197 101147 64225 101175
rect 64259 101147 64287 101175
rect 64321 101147 64349 101175
rect 64383 101147 64411 101175
rect 64197 101085 64225 101113
rect 64259 101085 64287 101113
rect 64321 101085 64349 101113
rect 64383 101085 64411 101113
rect 64197 101023 64225 101051
rect 64259 101023 64287 101051
rect 64321 101023 64349 101051
rect 64383 101023 64411 101051
rect 64197 100961 64225 100989
rect 64259 100961 64287 100989
rect 64321 100961 64349 100989
rect 64383 100961 64411 100989
rect 50697 95147 50725 95175
rect 50759 95147 50787 95175
rect 50821 95147 50849 95175
rect 50883 95147 50911 95175
rect 50697 95085 50725 95113
rect 50759 95085 50787 95113
rect 50821 95085 50849 95113
rect 50883 95085 50911 95113
rect 50697 95023 50725 95051
rect 50759 95023 50787 95051
rect 50821 95023 50849 95051
rect 50883 95023 50911 95051
rect 50697 94961 50725 94989
rect 50759 94961 50787 94989
rect 50821 94961 50849 94989
rect 50883 94961 50911 94989
rect 54659 95147 54687 95175
rect 54721 95147 54749 95175
rect 54659 95085 54687 95113
rect 54721 95085 54749 95113
rect 54659 95023 54687 95051
rect 54721 95023 54749 95051
rect 54659 94961 54687 94989
rect 54721 94961 54749 94989
rect 62339 92147 62367 92175
rect 62401 92147 62429 92175
rect 62339 92085 62367 92113
rect 62401 92085 62429 92113
rect 62339 92023 62367 92051
rect 62401 92023 62429 92051
rect 62339 91961 62367 91989
rect 62401 91961 62429 91989
rect 64197 92147 64225 92175
rect 64259 92147 64287 92175
rect 64321 92147 64349 92175
rect 64383 92147 64411 92175
rect 64197 92085 64225 92113
rect 64259 92085 64287 92113
rect 64321 92085 64349 92113
rect 64383 92085 64411 92113
rect 64197 92023 64225 92051
rect 64259 92023 64287 92051
rect 64321 92023 64349 92051
rect 64383 92023 64411 92051
rect 64197 91961 64225 91989
rect 64259 91961 64287 91989
rect 64321 91961 64349 91989
rect 64383 91961 64411 91989
rect 66057 167147 66085 167175
rect 66119 167147 66147 167175
rect 66181 167147 66209 167175
rect 66243 167147 66271 167175
rect 66057 167085 66085 167113
rect 66119 167085 66147 167113
rect 66181 167085 66209 167113
rect 66243 167085 66271 167113
rect 66057 167023 66085 167051
rect 66119 167023 66147 167051
rect 66181 167023 66209 167051
rect 66243 167023 66271 167051
rect 66057 166961 66085 166989
rect 66119 166961 66147 166989
rect 66181 166961 66209 166989
rect 66243 166961 66271 166989
rect 79557 164147 79585 164175
rect 79619 164147 79647 164175
rect 79681 164147 79709 164175
rect 79743 164147 79771 164175
rect 79557 164085 79585 164113
rect 79619 164085 79647 164113
rect 79681 164085 79709 164113
rect 79743 164085 79771 164113
rect 79557 164023 79585 164051
rect 79619 164023 79647 164051
rect 79681 164023 79709 164051
rect 79743 164023 79771 164051
rect 79557 163961 79585 163989
rect 79619 163961 79647 163989
rect 79681 163961 79709 163989
rect 79743 163961 79771 163989
rect 66057 158147 66085 158175
rect 66119 158147 66147 158175
rect 66181 158147 66209 158175
rect 66243 158147 66271 158175
rect 66057 158085 66085 158113
rect 66119 158085 66147 158113
rect 66181 158085 66209 158113
rect 66243 158085 66271 158113
rect 66057 158023 66085 158051
rect 66119 158023 66147 158051
rect 66181 158023 66209 158051
rect 66243 158023 66271 158051
rect 66057 157961 66085 157989
rect 66119 157961 66147 157989
rect 66181 157961 66209 157989
rect 66243 157961 66271 157989
rect 70659 158147 70687 158175
rect 70721 158147 70749 158175
rect 70659 158085 70687 158113
rect 70721 158085 70749 158113
rect 70659 158023 70687 158051
rect 70721 158023 70749 158051
rect 70659 157961 70687 157989
rect 70721 157961 70749 157989
rect 78339 155147 78367 155175
rect 78401 155147 78429 155175
rect 78339 155085 78367 155113
rect 78401 155085 78429 155113
rect 78339 155023 78367 155051
rect 78401 155023 78429 155051
rect 78339 154961 78367 154989
rect 78401 154961 78429 154989
rect 79557 155147 79585 155175
rect 79619 155147 79647 155175
rect 79681 155147 79709 155175
rect 79743 155147 79771 155175
rect 79557 155085 79585 155113
rect 79619 155085 79647 155113
rect 79681 155085 79709 155113
rect 79743 155085 79771 155113
rect 79557 155023 79585 155051
rect 79619 155023 79647 155051
rect 79681 155023 79709 155051
rect 79743 155023 79771 155051
rect 79557 154961 79585 154989
rect 79619 154961 79647 154989
rect 79681 154961 79709 154989
rect 79743 154961 79771 154989
rect 66057 149147 66085 149175
rect 66119 149147 66147 149175
rect 66181 149147 66209 149175
rect 66243 149147 66271 149175
rect 66057 149085 66085 149113
rect 66119 149085 66147 149113
rect 66181 149085 66209 149113
rect 66243 149085 66271 149113
rect 66057 149023 66085 149051
rect 66119 149023 66147 149051
rect 66181 149023 66209 149051
rect 66243 149023 66271 149051
rect 66057 148961 66085 148989
rect 66119 148961 66147 148989
rect 66181 148961 66209 148989
rect 66243 148961 66271 148989
rect 70659 149147 70687 149175
rect 70721 149147 70749 149175
rect 70659 149085 70687 149113
rect 70721 149085 70749 149113
rect 70659 149023 70687 149051
rect 70721 149023 70749 149051
rect 70659 148961 70687 148989
rect 70721 148961 70749 148989
rect 78339 146147 78367 146175
rect 78401 146147 78429 146175
rect 78339 146085 78367 146113
rect 78401 146085 78429 146113
rect 78339 146023 78367 146051
rect 78401 146023 78429 146051
rect 78339 145961 78367 145989
rect 78401 145961 78429 145989
rect 79557 146147 79585 146175
rect 79619 146147 79647 146175
rect 79681 146147 79709 146175
rect 79743 146147 79771 146175
rect 79557 146085 79585 146113
rect 79619 146085 79647 146113
rect 79681 146085 79709 146113
rect 79743 146085 79771 146113
rect 79557 146023 79585 146051
rect 79619 146023 79647 146051
rect 79681 146023 79709 146051
rect 79743 146023 79771 146051
rect 79557 145961 79585 145989
rect 79619 145961 79647 145989
rect 79681 145961 79709 145989
rect 79743 145961 79771 145989
rect 66057 140147 66085 140175
rect 66119 140147 66147 140175
rect 66181 140147 66209 140175
rect 66243 140147 66271 140175
rect 66057 140085 66085 140113
rect 66119 140085 66147 140113
rect 66181 140085 66209 140113
rect 66243 140085 66271 140113
rect 66057 140023 66085 140051
rect 66119 140023 66147 140051
rect 66181 140023 66209 140051
rect 66243 140023 66271 140051
rect 66057 139961 66085 139989
rect 66119 139961 66147 139989
rect 66181 139961 66209 139989
rect 66243 139961 66271 139989
rect 70659 140147 70687 140175
rect 70721 140147 70749 140175
rect 70659 140085 70687 140113
rect 70721 140085 70749 140113
rect 70659 140023 70687 140051
rect 70721 140023 70749 140051
rect 70659 139961 70687 139989
rect 70721 139961 70749 139989
rect 78339 137147 78367 137175
rect 78401 137147 78429 137175
rect 78339 137085 78367 137113
rect 78401 137085 78429 137113
rect 78339 137023 78367 137051
rect 78401 137023 78429 137051
rect 78339 136961 78367 136989
rect 78401 136961 78429 136989
rect 79557 137147 79585 137175
rect 79619 137147 79647 137175
rect 79681 137147 79709 137175
rect 79743 137147 79771 137175
rect 79557 137085 79585 137113
rect 79619 137085 79647 137113
rect 79681 137085 79709 137113
rect 79743 137085 79771 137113
rect 79557 137023 79585 137051
rect 79619 137023 79647 137051
rect 79681 137023 79709 137051
rect 79743 137023 79771 137051
rect 79557 136961 79585 136989
rect 79619 136961 79647 136989
rect 79681 136961 79709 136989
rect 79743 136961 79771 136989
rect 66057 131147 66085 131175
rect 66119 131147 66147 131175
rect 66181 131147 66209 131175
rect 66243 131147 66271 131175
rect 66057 131085 66085 131113
rect 66119 131085 66147 131113
rect 66181 131085 66209 131113
rect 66243 131085 66271 131113
rect 66057 131023 66085 131051
rect 66119 131023 66147 131051
rect 66181 131023 66209 131051
rect 66243 131023 66271 131051
rect 66057 130961 66085 130989
rect 66119 130961 66147 130989
rect 66181 130961 66209 130989
rect 66243 130961 66271 130989
rect 66057 122147 66085 122175
rect 66119 122147 66147 122175
rect 66181 122147 66209 122175
rect 66243 122147 66271 122175
rect 66057 122085 66085 122113
rect 66119 122085 66147 122113
rect 66181 122085 66209 122113
rect 66243 122085 66271 122113
rect 66057 122023 66085 122051
rect 66119 122023 66147 122051
rect 66181 122023 66209 122051
rect 66243 122023 66271 122051
rect 66057 121961 66085 121989
rect 66119 121961 66147 121989
rect 66181 121961 66209 121989
rect 66243 121961 66271 121989
rect 66057 113147 66085 113175
rect 66119 113147 66147 113175
rect 66181 113147 66209 113175
rect 66243 113147 66271 113175
rect 66057 113085 66085 113113
rect 66119 113085 66147 113113
rect 66181 113085 66209 113113
rect 66243 113085 66271 113113
rect 66057 113023 66085 113051
rect 66119 113023 66147 113051
rect 66181 113023 66209 113051
rect 66243 113023 66271 113051
rect 66057 112961 66085 112989
rect 66119 112961 66147 112989
rect 66181 112961 66209 112989
rect 66243 112961 66271 112989
rect 66057 104147 66085 104175
rect 66119 104147 66147 104175
rect 66181 104147 66209 104175
rect 66243 104147 66271 104175
rect 66057 104085 66085 104113
rect 66119 104085 66147 104113
rect 66181 104085 66209 104113
rect 66243 104085 66271 104113
rect 66057 104023 66085 104051
rect 66119 104023 66147 104051
rect 66181 104023 66209 104051
rect 66243 104023 66271 104051
rect 66057 103961 66085 103989
rect 66119 103961 66147 103989
rect 66181 103961 66209 103989
rect 66243 103961 66271 103989
rect 79557 128147 79585 128175
rect 79619 128147 79647 128175
rect 79681 128147 79709 128175
rect 79743 128147 79771 128175
rect 79557 128085 79585 128113
rect 79619 128085 79647 128113
rect 79681 128085 79709 128113
rect 79743 128085 79771 128113
rect 79557 128023 79585 128051
rect 79619 128023 79647 128051
rect 79681 128023 79709 128051
rect 79743 128023 79771 128051
rect 79557 127961 79585 127989
rect 79619 127961 79647 127989
rect 79681 127961 79709 127989
rect 79743 127961 79771 127989
rect 79557 119147 79585 119175
rect 79619 119147 79647 119175
rect 79681 119147 79709 119175
rect 79743 119147 79771 119175
rect 79557 119085 79585 119113
rect 79619 119085 79647 119113
rect 79681 119085 79709 119113
rect 79743 119085 79771 119113
rect 79557 119023 79585 119051
rect 79619 119023 79647 119051
rect 79681 119023 79709 119051
rect 79743 119023 79771 119051
rect 79557 118961 79585 118989
rect 79619 118961 79647 118989
rect 79681 118961 79709 118989
rect 79743 118961 79771 118989
rect 79557 110147 79585 110175
rect 79619 110147 79647 110175
rect 79681 110147 79709 110175
rect 79743 110147 79771 110175
rect 79557 110085 79585 110113
rect 79619 110085 79647 110113
rect 79681 110085 79709 110113
rect 79743 110085 79771 110113
rect 79557 110023 79585 110051
rect 79619 110023 79647 110051
rect 79681 110023 79709 110051
rect 79743 110023 79771 110051
rect 79557 109961 79585 109989
rect 79619 109961 79647 109989
rect 79681 109961 79709 109989
rect 79743 109961 79771 109989
rect 77699 101147 77727 101175
rect 77761 101147 77789 101175
rect 77699 101085 77727 101113
rect 77761 101085 77789 101113
rect 77699 101023 77727 101051
rect 77761 101023 77789 101051
rect 77699 100961 77727 100989
rect 77761 100961 77789 100989
rect 79557 101147 79585 101175
rect 79619 101147 79647 101175
rect 79681 101147 79709 101175
rect 79743 101147 79771 101175
rect 79557 101085 79585 101113
rect 79619 101085 79647 101113
rect 79681 101085 79709 101113
rect 79743 101085 79771 101113
rect 79557 101023 79585 101051
rect 79619 101023 79647 101051
rect 79681 101023 79709 101051
rect 79743 101023 79771 101051
rect 79557 100961 79585 100989
rect 79619 100961 79647 100989
rect 79681 100961 79709 100989
rect 79743 100961 79771 100989
rect 66057 95147 66085 95175
rect 66119 95147 66147 95175
rect 66181 95147 66209 95175
rect 66243 95147 66271 95175
rect 66057 95085 66085 95113
rect 66119 95085 66147 95113
rect 66181 95085 66209 95113
rect 66243 95085 66271 95113
rect 66057 95023 66085 95051
rect 66119 95023 66147 95051
rect 66181 95023 66209 95051
rect 66243 95023 66271 95051
rect 66057 94961 66085 94989
rect 66119 94961 66147 94989
rect 66181 94961 66209 94989
rect 66243 94961 66271 94989
rect 70019 95147 70047 95175
rect 70081 95147 70109 95175
rect 70019 95085 70047 95113
rect 70081 95085 70109 95113
rect 70019 95023 70047 95051
rect 70081 95023 70109 95051
rect 70019 94961 70047 94989
rect 70081 94961 70109 94989
rect 77699 92147 77727 92175
rect 77761 92147 77789 92175
rect 77699 92085 77727 92113
rect 77761 92085 77789 92113
rect 77699 92023 77727 92051
rect 77761 92023 77789 92051
rect 77699 91961 77727 91989
rect 77761 91961 77789 91989
rect 79557 92147 79585 92175
rect 79619 92147 79647 92175
rect 79681 92147 79709 92175
rect 79743 92147 79771 92175
rect 79557 92085 79585 92113
rect 79619 92085 79647 92113
rect 79681 92085 79709 92113
rect 79743 92085 79771 92113
rect 79557 92023 79585 92051
rect 79619 92023 79647 92051
rect 79681 92023 79709 92051
rect 79743 92023 79771 92051
rect 79557 91961 79585 91989
rect 79619 91961 79647 91989
rect 79681 91961 79709 91989
rect 79743 91961 79771 91989
rect 23939 86147 23967 86175
rect 24001 86147 24029 86175
rect 23939 86085 23967 86113
rect 24001 86085 24029 86113
rect 23939 86023 23967 86051
rect 24001 86023 24029 86051
rect 23939 85961 23967 85989
rect 24001 85961 24029 85989
rect 39299 86147 39327 86175
rect 39361 86147 39389 86175
rect 39299 86085 39327 86113
rect 39361 86085 39389 86113
rect 39299 86023 39327 86051
rect 39361 86023 39389 86051
rect 39299 85961 39327 85989
rect 39361 85961 39389 85989
rect 54659 86147 54687 86175
rect 54721 86147 54749 86175
rect 54659 86085 54687 86113
rect 54721 86085 54749 86113
rect 54659 86023 54687 86051
rect 54721 86023 54749 86051
rect 54659 85961 54687 85989
rect 54721 85961 54749 85989
rect 70019 86147 70047 86175
rect 70081 86147 70109 86175
rect 70019 86085 70047 86113
rect 70081 86085 70109 86113
rect 70019 86023 70047 86051
rect 70081 86023 70109 86051
rect 70019 85961 70047 85989
rect 70081 85961 70109 85989
rect 31619 83147 31647 83175
rect 31681 83147 31709 83175
rect 31619 83085 31647 83113
rect 31681 83085 31709 83113
rect 31619 83023 31647 83051
rect 31681 83023 31709 83051
rect 31619 82961 31647 82989
rect 31681 82961 31709 82989
rect 46979 83147 47007 83175
rect 47041 83147 47069 83175
rect 46979 83085 47007 83113
rect 47041 83085 47069 83113
rect 46979 83023 47007 83051
rect 47041 83023 47069 83051
rect 46979 82961 47007 82989
rect 47041 82961 47069 82989
rect 62339 83147 62367 83175
rect 62401 83147 62429 83175
rect 62339 83085 62367 83113
rect 62401 83085 62429 83113
rect 62339 83023 62367 83051
rect 62401 83023 62429 83051
rect 62339 82961 62367 82989
rect 62401 82961 62429 82989
rect 77699 83147 77727 83175
rect 77761 83147 77789 83175
rect 77699 83085 77727 83113
rect 77761 83085 77789 83113
rect 77699 83023 77727 83051
rect 77761 83023 77789 83051
rect 77699 82961 77727 82989
rect 77761 82961 77789 82989
rect 79557 83147 79585 83175
rect 79619 83147 79647 83175
rect 79681 83147 79709 83175
rect 79743 83147 79771 83175
rect 79557 83085 79585 83113
rect 79619 83085 79647 83113
rect 79681 83085 79709 83113
rect 79743 83085 79771 83113
rect 79557 83023 79585 83051
rect 79619 83023 79647 83051
rect 79681 83023 79709 83051
rect 79743 83023 79771 83051
rect 79557 82961 79585 82989
rect 79619 82961 79647 82989
rect 79681 82961 79709 82989
rect 79743 82961 79771 82989
rect 23939 77147 23967 77175
rect 24001 77147 24029 77175
rect 23939 77085 23967 77113
rect 24001 77085 24029 77113
rect 23939 77023 23967 77051
rect 24001 77023 24029 77051
rect 23939 76961 23967 76989
rect 24001 76961 24029 76989
rect 39299 77147 39327 77175
rect 39361 77147 39389 77175
rect 39299 77085 39327 77113
rect 39361 77085 39389 77113
rect 39299 77023 39327 77051
rect 39361 77023 39389 77051
rect 39299 76961 39327 76989
rect 39361 76961 39389 76989
rect 54659 77147 54687 77175
rect 54721 77147 54749 77175
rect 54659 77085 54687 77113
rect 54721 77085 54749 77113
rect 54659 77023 54687 77051
rect 54721 77023 54749 77051
rect 54659 76961 54687 76989
rect 54721 76961 54749 76989
rect 70019 77147 70047 77175
rect 70081 77147 70109 77175
rect 70019 77085 70047 77113
rect 70081 77085 70109 77113
rect 70019 77023 70047 77051
rect 70081 77023 70109 77051
rect 70019 76961 70047 76989
rect 70081 76961 70109 76989
rect 19977 68147 20005 68175
rect 20039 68147 20067 68175
rect 20101 68147 20129 68175
rect 20163 68147 20191 68175
rect 19977 68085 20005 68113
rect 20039 68085 20067 68113
rect 20101 68085 20129 68113
rect 20163 68085 20191 68113
rect 19977 68023 20005 68051
rect 20039 68023 20067 68051
rect 20101 68023 20129 68051
rect 20163 68023 20191 68051
rect 19977 67961 20005 67989
rect 20039 67961 20067 67989
rect 20101 67961 20129 67989
rect 20163 67961 20191 67989
rect 19977 59147 20005 59175
rect 20039 59147 20067 59175
rect 20101 59147 20129 59175
rect 20163 59147 20191 59175
rect 19977 59085 20005 59113
rect 20039 59085 20067 59113
rect 20101 59085 20129 59113
rect 20163 59085 20191 59113
rect 19977 59023 20005 59051
rect 20039 59023 20067 59051
rect 20101 59023 20129 59051
rect 20163 59023 20191 59051
rect 19977 58961 20005 58989
rect 20039 58961 20067 58989
rect 20101 58961 20129 58989
rect 20163 58961 20191 58989
rect 19977 50147 20005 50175
rect 20039 50147 20067 50175
rect 20101 50147 20129 50175
rect 20163 50147 20191 50175
rect 19977 50085 20005 50113
rect 20039 50085 20067 50113
rect 20101 50085 20129 50113
rect 20163 50085 20191 50113
rect 19977 50023 20005 50051
rect 20039 50023 20067 50051
rect 20101 50023 20129 50051
rect 20163 50023 20191 50051
rect 19977 49961 20005 49989
rect 20039 49961 20067 49989
rect 20101 49961 20129 49989
rect 20163 49961 20191 49989
rect 19977 41147 20005 41175
rect 20039 41147 20067 41175
rect 20101 41147 20129 41175
rect 20163 41147 20191 41175
rect 19977 41085 20005 41113
rect 20039 41085 20067 41113
rect 20101 41085 20129 41113
rect 20163 41085 20191 41113
rect 19977 41023 20005 41051
rect 20039 41023 20067 41051
rect 20101 41023 20129 41051
rect 20163 41023 20191 41051
rect 19977 40961 20005 40989
rect 20039 40961 20067 40989
rect 20101 40961 20129 40989
rect 20163 40961 20191 40989
rect 19977 32147 20005 32175
rect 20039 32147 20067 32175
rect 20101 32147 20129 32175
rect 20163 32147 20191 32175
rect 19977 32085 20005 32113
rect 20039 32085 20067 32113
rect 20101 32085 20129 32113
rect 20163 32085 20191 32113
rect 19977 32023 20005 32051
rect 20039 32023 20067 32051
rect 20101 32023 20129 32051
rect 20163 32023 20191 32051
rect 19977 31961 20005 31989
rect 20039 31961 20067 31989
rect 20101 31961 20129 31989
rect 20163 31961 20191 31989
rect 19977 23147 20005 23175
rect 20039 23147 20067 23175
rect 20101 23147 20129 23175
rect 20163 23147 20191 23175
rect 19977 23085 20005 23113
rect 20039 23085 20067 23113
rect 20101 23085 20129 23113
rect 20163 23085 20191 23113
rect 19977 23023 20005 23051
rect 20039 23023 20067 23051
rect 20101 23023 20129 23051
rect 20163 23023 20191 23051
rect 19977 22961 20005 22989
rect 20039 22961 20067 22989
rect 20101 22961 20129 22989
rect 20163 22961 20191 22989
rect 19977 14147 20005 14175
rect 20039 14147 20067 14175
rect 20101 14147 20129 14175
rect 20163 14147 20191 14175
rect 19977 14085 20005 14113
rect 20039 14085 20067 14113
rect 20101 14085 20129 14113
rect 20163 14085 20191 14113
rect 19977 14023 20005 14051
rect 20039 14023 20067 14051
rect 20101 14023 20129 14051
rect 20163 14023 20191 14051
rect 19977 13961 20005 13989
rect 20039 13961 20067 13989
rect 20101 13961 20129 13989
rect 20163 13961 20191 13989
rect 19977 5147 20005 5175
rect 20039 5147 20067 5175
rect 20101 5147 20129 5175
rect 20163 5147 20191 5175
rect 19977 5085 20005 5113
rect 20039 5085 20067 5113
rect 20101 5085 20129 5113
rect 20163 5085 20191 5113
rect 19977 5023 20005 5051
rect 20039 5023 20067 5051
rect 20101 5023 20129 5051
rect 20163 5023 20191 5051
rect 19977 4961 20005 4989
rect 20039 4961 20067 4989
rect 20101 4961 20129 4989
rect 20163 4961 20191 4989
rect 19977 -588 20005 -560
rect 20039 -588 20067 -560
rect 20101 -588 20129 -560
rect 20163 -588 20191 -560
rect 19977 -650 20005 -622
rect 20039 -650 20067 -622
rect 20101 -650 20129 -622
rect 20163 -650 20191 -622
rect 19977 -712 20005 -684
rect 20039 -712 20067 -684
rect 20101 -712 20129 -684
rect 20163 -712 20191 -684
rect 19977 -774 20005 -746
rect 20039 -774 20067 -746
rect 20101 -774 20129 -746
rect 20163 -774 20191 -746
rect 33477 74147 33505 74175
rect 33539 74147 33567 74175
rect 33601 74147 33629 74175
rect 33663 74147 33691 74175
rect 33477 74085 33505 74113
rect 33539 74085 33567 74113
rect 33601 74085 33629 74113
rect 33663 74085 33691 74113
rect 33477 74023 33505 74051
rect 33539 74023 33567 74051
rect 33601 74023 33629 74051
rect 33663 74023 33691 74051
rect 33477 73961 33505 73989
rect 33539 73961 33567 73989
rect 33601 73961 33629 73989
rect 33663 73961 33691 73989
rect 33477 65147 33505 65175
rect 33539 65147 33567 65175
rect 33601 65147 33629 65175
rect 33663 65147 33691 65175
rect 33477 65085 33505 65113
rect 33539 65085 33567 65113
rect 33601 65085 33629 65113
rect 33663 65085 33691 65113
rect 33477 65023 33505 65051
rect 33539 65023 33567 65051
rect 33601 65023 33629 65051
rect 33663 65023 33691 65051
rect 33477 64961 33505 64989
rect 33539 64961 33567 64989
rect 33601 64961 33629 64989
rect 33663 64961 33691 64989
rect 33477 56147 33505 56175
rect 33539 56147 33567 56175
rect 33601 56147 33629 56175
rect 33663 56147 33691 56175
rect 33477 56085 33505 56113
rect 33539 56085 33567 56113
rect 33601 56085 33629 56113
rect 33663 56085 33691 56113
rect 33477 56023 33505 56051
rect 33539 56023 33567 56051
rect 33601 56023 33629 56051
rect 33663 56023 33691 56051
rect 33477 55961 33505 55989
rect 33539 55961 33567 55989
rect 33601 55961 33629 55989
rect 33663 55961 33691 55989
rect 33477 47147 33505 47175
rect 33539 47147 33567 47175
rect 33601 47147 33629 47175
rect 33663 47147 33691 47175
rect 33477 47085 33505 47113
rect 33539 47085 33567 47113
rect 33601 47085 33629 47113
rect 33663 47085 33691 47113
rect 33477 47023 33505 47051
rect 33539 47023 33567 47051
rect 33601 47023 33629 47051
rect 33663 47023 33691 47051
rect 33477 46961 33505 46989
rect 33539 46961 33567 46989
rect 33601 46961 33629 46989
rect 33663 46961 33691 46989
rect 33477 38147 33505 38175
rect 33539 38147 33567 38175
rect 33601 38147 33629 38175
rect 33663 38147 33691 38175
rect 33477 38085 33505 38113
rect 33539 38085 33567 38113
rect 33601 38085 33629 38113
rect 33663 38085 33691 38113
rect 33477 38023 33505 38051
rect 33539 38023 33567 38051
rect 33601 38023 33629 38051
rect 33663 38023 33691 38051
rect 33477 37961 33505 37989
rect 33539 37961 33567 37989
rect 33601 37961 33629 37989
rect 33663 37961 33691 37989
rect 33477 29147 33505 29175
rect 33539 29147 33567 29175
rect 33601 29147 33629 29175
rect 33663 29147 33691 29175
rect 33477 29085 33505 29113
rect 33539 29085 33567 29113
rect 33601 29085 33629 29113
rect 33663 29085 33691 29113
rect 33477 29023 33505 29051
rect 33539 29023 33567 29051
rect 33601 29023 33629 29051
rect 33663 29023 33691 29051
rect 33477 28961 33505 28989
rect 33539 28961 33567 28989
rect 33601 28961 33629 28989
rect 33663 28961 33691 28989
rect 33477 20147 33505 20175
rect 33539 20147 33567 20175
rect 33601 20147 33629 20175
rect 33663 20147 33691 20175
rect 33477 20085 33505 20113
rect 33539 20085 33567 20113
rect 33601 20085 33629 20113
rect 33663 20085 33691 20113
rect 33477 20023 33505 20051
rect 33539 20023 33567 20051
rect 33601 20023 33629 20051
rect 33663 20023 33691 20051
rect 33477 19961 33505 19989
rect 33539 19961 33567 19989
rect 33601 19961 33629 19989
rect 33663 19961 33691 19989
rect 33477 11147 33505 11175
rect 33539 11147 33567 11175
rect 33601 11147 33629 11175
rect 33663 11147 33691 11175
rect 33477 11085 33505 11113
rect 33539 11085 33567 11113
rect 33601 11085 33629 11113
rect 33663 11085 33691 11113
rect 33477 11023 33505 11051
rect 33539 11023 33567 11051
rect 33601 11023 33629 11051
rect 33663 11023 33691 11051
rect 33477 10961 33505 10989
rect 33539 10961 33567 10989
rect 33601 10961 33629 10989
rect 33663 10961 33691 10989
rect 33477 2147 33505 2175
rect 33539 2147 33567 2175
rect 33601 2147 33629 2175
rect 33663 2147 33691 2175
rect 33477 2085 33505 2113
rect 33539 2085 33567 2113
rect 33601 2085 33629 2113
rect 33663 2085 33691 2113
rect 33477 2023 33505 2051
rect 33539 2023 33567 2051
rect 33601 2023 33629 2051
rect 33663 2023 33691 2051
rect 33477 1961 33505 1989
rect 33539 1961 33567 1989
rect 33601 1961 33629 1989
rect 33663 1961 33691 1989
rect 33477 -108 33505 -80
rect 33539 -108 33567 -80
rect 33601 -108 33629 -80
rect 33663 -108 33691 -80
rect 33477 -170 33505 -142
rect 33539 -170 33567 -142
rect 33601 -170 33629 -142
rect 33663 -170 33691 -142
rect 33477 -232 33505 -204
rect 33539 -232 33567 -204
rect 33601 -232 33629 -204
rect 33663 -232 33691 -204
rect 33477 -294 33505 -266
rect 33539 -294 33567 -266
rect 33601 -294 33629 -266
rect 33663 -294 33691 -266
rect 35337 68147 35365 68175
rect 35399 68147 35427 68175
rect 35461 68147 35489 68175
rect 35523 68147 35551 68175
rect 35337 68085 35365 68113
rect 35399 68085 35427 68113
rect 35461 68085 35489 68113
rect 35523 68085 35551 68113
rect 35337 68023 35365 68051
rect 35399 68023 35427 68051
rect 35461 68023 35489 68051
rect 35523 68023 35551 68051
rect 35337 67961 35365 67989
rect 35399 67961 35427 67989
rect 35461 67961 35489 67989
rect 35523 67961 35551 67989
rect 35337 59147 35365 59175
rect 35399 59147 35427 59175
rect 35461 59147 35489 59175
rect 35523 59147 35551 59175
rect 35337 59085 35365 59113
rect 35399 59085 35427 59113
rect 35461 59085 35489 59113
rect 35523 59085 35551 59113
rect 35337 59023 35365 59051
rect 35399 59023 35427 59051
rect 35461 59023 35489 59051
rect 35523 59023 35551 59051
rect 35337 58961 35365 58989
rect 35399 58961 35427 58989
rect 35461 58961 35489 58989
rect 35523 58961 35551 58989
rect 35337 50147 35365 50175
rect 35399 50147 35427 50175
rect 35461 50147 35489 50175
rect 35523 50147 35551 50175
rect 35337 50085 35365 50113
rect 35399 50085 35427 50113
rect 35461 50085 35489 50113
rect 35523 50085 35551 50113
rect 35337 50023 35365 50051
rect 35399 50023 35427 50051
rect 35461 50023 35489 50051
rect 35523 50023 35551 50051
rect 35337 49961 35365 49989
rect 35399 49961 35427 49989
rect 35461 49961 35489 49989
rect 35523 49961 35551 49989
rect 35337 41147 35365 41175
rect 35399 41147 35427 41175
rect 35461 41147 35489 41175
rect 35523 41147 35551 41175
rect 35337 41085 35365 41113
rect 35399 41085 35427 41113
rect 35461 41085 35489 41113
rect 35523 41085 35551 41113
rect 35337 41023 35365 41051
rect 35399 41023 35427 41051
rect 35461 41023 35489 41051
rect 35523 41023 35551 41051
rect 35337 40961 35365 40989
rect 35399 40961 35427 40989
rect 35461 40961 35489 40989
rect 35523 40961 35551 40989
rect 35337 32147 35365 32175
rect 35399 32147 35427 32175
rect 35461 32147 35489 32175
rect 35523 32147 35551 32175
rect 35337 32085 35365 32113
rect 35399 32085 35427 32113
rect 35461 32085 35489 32113
rect 35523 32085 35551 32113
rect 35337 32023 35365 32051
rect 35399 32023 35427 32051
rect 35461 32023 35489 32051
rect 35523 32023 35551 32051
rect 35337 31961 35365 31989
rect 35399 31961 35427 31989
rect 35461 31961 35489 31989
rect 35523 31961 35551 31989
rect 35337 23147 35365 23175
rect 35399 23147 35427 23175
rect 35461 23147 35489 23175
rect 35523 23147 35551 23175
rect 35337 23085 35365 23113
rect 35399 23085 35427 23113
rect 35461 23085 35489 23113
rect 35523 23085 35551 23113
rect 35337 23023 35365 23051
rect 35399 23023 35427 23051
rect 35461 23023 35489 23051
rect 35523 23023 35551 23051
rect 35337 22961 35365 22989
rect 35399 22961 35427 22989
rect 35461 22961 35489 22989
rect 35523 22961 35551 22989
rect 35337 14147 35365 14175
rect 35399 14147 35427 14175
rect 35461 14147 35489 14175
rect 35523 14147 35551 14175
rect 35337 14085 35365 14113
rect 35399 14085 35427 14113
rect 35461 14085 35489 14113
rect 35523 14085 35551 14113
rect 35337 14023 35365 14051
rect 35399 14023 35427 14051
rect 35461 14023 35489 14051
rect 35523 14023 35551 14051
rect 35337 13961 35365 13989
rect 35399 13961 35427 13989
rect 35461 13961 35489 13989
rect 35523 13961 35551 13989
rect 35337 5147 35365 5175
rect 35399 5147 35427 5175
rect 35461 5147 35489 5175
rect 35523 5147 35551 5175
rect 35337 5085 35365 5113
rect 35399 5085 35427 5113
rect 35461 5085 35489 5113
rect 35523 5085 35551 5113
rect 35337 5023 35365 5051
rect 35399 5023 35427 5051
rect 35461 5023 35489 5051
rect 35523 5023 35551 5051
rect 35337 4961 35365 4989
rect 35399 4961 35427 4989
rect 35461 4961 35489 4989
rect 35523 4961 35551 4989
rect 35337 -588 35365 -560
rect 35399 -588 35427 -560
rect 35461 -588 35489 -560
rect 35523 -588 35551 -560
rect 35337 -650 35365 -622
rect 35399 -650 35427 -622
rect 35461 -650 35489 -622
rect 35523 -650 35551 -622
rect 35337 -712 35365 -684
rect 35399 -712 35427 -684
rect 35461 -712 35489 -684
rect 35523 -712 35551 -684
rect 35337 -774 35365 -746
rect 35399 -774 35427 -746
rect 35461 -774 35489 -746
rect 35523 -774 35551 -746
rect 48837 74147 48865 74175
rect 48899 74147 48927 74175
rect 48961 74147 48989 74175
rect 49023 74147 49051 74175
rect 48837 74085 48865 74113
rect 48899 74085 48927 74113
rect 48961 74085 48989 74113
rect 49023 74085 49051 74113
rect 48837 74023 48865 74051
rect 48899 74023 48927 74051
rect 48961 74023 48989 74051
rect 49023 74023 49051 74051
rect 48837 73961 48865 73989
rect 48899 73961 48927 73989
rect 48961 73961 48989 73989
rect 49023 73961 49051 73989
rect 48837 65147 48865 65175
rect 48899 65147 48927 65175
rect 48961 65147 48989 65175
rect 49023 65147 49051 65175
rect 48837 65085 48865 65113
rect 48899 65085 48927 65113
rect 48961 65085 48989 65113
rect 49023 65085 49051 65113
rect 48837 65023 48865 65051
rect 48899 65023 48927 65051
rect 48961 65023 48989 65051
rect 49023 65023 49051 65051
rect 48837 64961 48865 64989
rect 48899 64961 48927 64989
rect 48961 64961 48989 64989
rect 49023 64961 49051 64989
rect 48837 56147 48865 56175
rect 48899 56147 48927 56175
rect 48961 56147 48989 56175
rect 49023 56147 49051 56175
rect 48837 56085 48865 56113
rect 48899 56085 48927 56113
rect 48961 56085 48989 56113
rect 49023 56085 49051 56113
rect 48837 56023 48865 56051
rect 48899 56023 48927 56051
rect 48961 56023 48989 56051
rect 49023 56023 49051 56051
rect 48837 55961 48865 55989
rect 48899 55961 48927 55989
rect 48961 55961 48989 55989
rect 49023 55961 49051 55989
rect 48837 47147 48865 47175
rect 48899 47147 48927 47175
rect 48961 47147 48989 47175
rect 49023 47147 49051 47175
rect 48837 47085 48865 47113
rect 48899 47085 48927 47113
rect 48961 47085 48989 47113
rect 49023 47085 49051 47113
rect 48837 47023 48865 47051
rect 48899 47023 48927 47051
rect 48961 47023 48989 47051
rect 49023 47023 49051 47051
rect 48837 46961 48865 46989
rect 48899 46961 48927 46989
rect 48961 46961 48989 46989
rect 49023 46961 49051 46989
rect 48837 38147 48865 38175
rect 48899 38147 48927 38175
rect 48961 38147 48989 38175
rect 49023 38147 49051 38175
rect 48837 38085 48865 38113
rect 48899 38085 48927 38113
rect 48961 38085 48989 38113
rect 49023 38085 49051 38113
rect 48837 38023 48865 38051
rect 48899 38023 48927 38051
rect 48961 38023 48989 38051
rect 49023 38023 49051 38051
rect 48837 37961 48865 37989
rect 48899 37961 48927 37989
rect 48961 37961 48989 37989
rect 49023 37961 49051 37989
rect 48837 29147 48865 29175
rect 48899 29147 48927 29175
rect 48961 29147 48989 29175
rect 49023 29147 49051 29175
rect 48837 29085 48865 29113
rect 48899 29085 48927 29113
rect 48961 29085 48989 29113
rect 49023 29085 49051 29113
rect 48837 29023 48865 29051
rect 48899 29023 48927 29051
rect 48961 29023 48989 29051
rect 49023 29023 49051 29051
rect 48837 28961 48865 28989
rect 48899 28961 48927 28989
rect 48961 28961 48989 28989
rect 49023 28961 49051 28989
rect 48837 20147 48865 20175
rect 48899 20147 48927 20175
rect 48961 20147 48989 20175
rect 49023 20147 49051 20175
rect 48837 20085 48865 20113
rect 48899 20085 48927 20113
rect 48961 20085 48989 20113
rect 49023 20085 49051 20113
rect 48837 20023 48865 20051
rect 48899 20023 48927 20051
rect 48961 20023 48989 20051
rect 49023 20023 49051 20051
rect 48837 19961 48865 19989
rect 48899 19961 48927 19989
rect 48961 19961 48989 19989
rect 49023 19961 49051 19989
rect 48837 11147 48865 11175
rect 48899 11147 48927 11175
rect 48961 11147 48989 11175
rect 49023 11147 49051 11175
rect 48837 11085 48865 11113
rect 48899 11085 48927 11113
rect 48961 11085 48989 11113
rect 49023 11085 49051 11113
rect 48837 11023 48865 11051
rect 48899 11023 48927 11051
rect 48961 11023 48989 11051
rect 49023 11023 49051 11051
rect 48837 10961 48865 10989
rect 48899 10961 48927 10989
rect 48961 10961 48989 10989
rect 49023 10961 49051 10989
rect 48837 2147 48865 2175
rect 48899 2147 48927 2175
rect 48961 2147 48989 2175
rect 49023 2147 49051 2175
rect 48837 2085 48865 2113
rect 48899 2085 48927 2113
rect 48961 2085 48989 2113
rect 49023 2085 49051 2113
rect 48837 2023 48865 2051
rect 48899 2023 48927 2051
rect 48961 2023 48989 2051
rect 49023 2023 49051 2051
rect 48837 1961 48865 1989
rect 48899 1961 48927 1989
rect 48961 1961 48989 1989
rect 49023 1961 49051 1989
rect 48837 -108 48865 -80
rect 48899 -108 48927 -80
rect 48961 -108 48989 -80
rect 49023 -108 49051 -80
rect 48837 -170 48865 -142
rect 48899 -170 48927 -142
rect 48961 -170 48989 -142
rect 49023 -170 49051 -142
rect 48837 -232 48865 -204
rect 48899 -232 48927 -204
rect 48961 -232 48989 -204
rect 49023 -232 49051 -204
rect 48837 -294 48865 -266
rect 48899 -294 48927 -266
rect 48961 -294 48989 -266
rect 49023 -294 49051 -266
rect 50697 68147 50725 68175
rect 50759 68147 50787 68175
rect 50821 68147 50849 68175
rect 50883 68147 50911 68175
rect 50697 68085 50725 68113
rect 50759 68085 50787 68113
rect 50821 68085 50849 68113
rect 50883 68085 50911 68113
rect 50697 68023 50725 68051
rect 50759 68023 50787 68051
rect 50821 68023 50849 68051
rect 50883 68023 50911 68051
rect 50697 67961 50725 67989
rect 50759 67961 50787 67989
rect 50821 67961 50849 67989
rect 50883 67961 50911 67989
rect 50697 59147 50725 59175
rect 50759 59147 50787 59175
rect 50821 59147 50849 59175
rect 50883 59147 50911 59175
rect 50697 59085 50725 59113
rect 50759 59085 50787 59113
rect 50821 59085 50849 59113
rect 50883 59085 50911 59113
rect 50697 59023 50725 59051
rect 50759 59023 50787 59051
rect 50821 59023 50849 59051
rect 50883 59023 50911 59051
rect 50697 58961 50725 58989
rect 50759 58961 50787 58989
rect 50821 58961 50849 58989
rect 50883 58961 50911 58989
rect 50697 50147 50725 50175
rect 50759 50147 50787 50175
rect 50821 50147 50849 50175
rect 50883 50147 50911 50175
rect 50697 50085 50725 50113
rect 50759 50085 50787 50113
rect 50821 50085 50849 50113
rect 50883 50085 50911 50113
rect 50697 50023 50725 50051
rect 50759 50023 50787 50051
rect 50821 50023 50849 50051
rect 50883 50023 50911 50051
rect 50697 49961 50725 49989
rect 50759 49961 50787 49989
rect 50821 49961 50849 49989
rect 50883 49961 50911 49989
rect 50697 41147 50725 41175
rect 50759 41147 50787 41175
rect 50821 41147 50849 41175
rect 50883 41147 50911 41175
rect 50697 41085 50725 41113
rect 50759 41085 50787 41113
rect 50821 41085 50849 41113
rect 50883 41085 50911 41113
rect 50697 41023 50725 41051
rect 50759 41023 50787 41051
rect 50821 41023 50849 41051
rect 50883 41023 50911 41051
rect 50697 40961 50725 40989
rect 50759 40961 50787 40989
rect 50821 40961 50849 40989
rect 50883 40961 50911 40989
rect 50697 32147 50725 32175
rect 50759 32147 50787 32175
rect 50821 32147 50849 32175
rect 50883 32147 50911 32175
rect 50697 32085 50725 32113
rect 50759 32085 50787 32113
rect 50821 32085 50849 32113
rect 50883 32085 50911 32113
rect 50697 32023 50725 32051
rect 50759 32023 50787 32051
rect 50821 32023 50849 32051
rect 50883 32023 50911 32051
rect 50697 31961 50725 31989
rect 50759 31961 50787 31989
rect 50821 31961 50849 31989
rect 50883 31961 50911 31989
rect 50697 23147 50725 23175
rect 50759 23147 50787 23175
rect 50821 23147 50849 23175
rect 50883 23147 50911 23175
rect 50697 23085 50725 23113
rect 50759 23085 50787 23113
rect 50821 23085 50849 23113
rect 50883 23085 50911 23113
rect 50697 23023 50725 23051
rect 50759 23023 50787 23051
rect 50821 23023 50849 23051
rect 50883 23023 50911 23051
rect 50697 22961 50725 22989
rect 50759 22961 50787 22989
rect 50821 22961 50849 22989
rect 50883 22961 50911 22989
rect 50697 14147 50725 14175
rect 50759 14147 50787 14175
rect 50821 14147 50849 14175
rect 50883 14147 50911 14175
rect 50697 14085 50725 14113
rect 50759 14085 50787 14113
rect 50821 14085 50849 14113
rect 50883 14085 50911 14113
rect 50697 14023 50725 14051
rect 50759 14023 50787 14051
rect 50821 14023 50849 14051
rect 50883 14023 50911 14051
rect 50697 13961 50725 13989
rect 50759 13961 50787 13989
rect 50821 13961 50849 13989
rect 50883 13961 50911 13989
rect 50697 5147 50725 5175
rect 50759 5147 50787 5175
rect 50821 5147 50849 5175
rect 50883 5147 50911 5175
rect 50697 5085 50725 5113
rect 50759 5085 50787 5113
rect 50821 5085 50849 5113
rect 50883 5085 50911 5113
rect 50697 5023 50725 5051
rect 50759 5023 50787 5051
rect 50821 5023 50849 5051
rect 50883 5023 50911 5051
rect 50697 4961 50725 4989
rect 50759 4961 50787 4989
rect 50821 4961 50849 4989
rect 50883 4961 50911 4989
rect 50697 -588 50725 -560
rect 50759 -588 50787 -560
rect 50821 -588 50849 -560
rect 50883 -588 50911 -560
rect 50697 -650 50725 -622
rect 50759 -650 50787 -622
rect 50821 -650 50849 -622
rect 50883 -650 50911 -622
rect 50697 -712 50725 -684
rect 50759 -712 50787 -684
rect 50821 -712 50849 -684
rect 50883 -712 50911 -684
rect 50697 -774 50725 -746
rect 50759 -774 50787 -746
rect 50821 -774 50849 -746
rect 50883 -774 50911 -746
rect 64197 74147 64225 74175
rect 64259 74147 64287 74175
rect 64321 74147 64349 74175
rect 64383 74147 64411 74175
rect 64197 74085 64225 74113
rect 64259 74085 64287 74113
rect 64321 74085 64349 74113
rect 64383 74085 64411 74113
rect 64197 74023 64225 74051
rect 64259 74023 64287 74051
rect 64321 74023 64349 74051
rect 64383 74023 64411 74051
rect 64197 73961 64225 73989
rect 64259 73961 64287 73989
rect 64321 73961 64349 73989
rect 64383 73961 64411 73989
rect 64197 65147 64225 65175
rect 64259 65147 64287 65175
rect 64321 65147 64349 65175
rect 64383 65147 64411 65175
rect 64197 65085 64225 65113
rect 64259 65085 64287 65113
rect 64321 65085 64349 65113
rect 64383 65085 64411 65113
rect 64197 65023 64225 65051
rect 64259 65023 64287 65051
rect 64321 65023 64349 65051
rect 64383 65023 64411 65051
rect 64197 64961 64225 64989
rect 64259 64961 64287 64989
rect 64321 64961 64349 64989
rect 64383 64961 64411 64989
rect 64197 56147 64225 56175
rect 64259 56147 64287 56175
rect 64321 56147 64349 56175
rect 64383 56147 64411 56175
rect 64197 56085 64225 56113
rect 64259 56085 64287 56113
rect 64321 56085 64349 56113
rect 64383 56085 64411 56113
rect 64197 56023 64225 56051
rect 64259 56023 64287 56051
rect 64321 56023 64349 56051
rect 64383 56023 64411 56051
rect 64197 55961 64225 55989
rect 64259 55961 64287 55989
rect 64321 55961 64349 55989
rect 64383 55961 64411 55989
rect 64197 47147 64225 47175
rect 64259 47147 64287 47175
rect 64321 47147 64349 47175
rect 64383 47147 64411 47175
rect 64197 47085 64225 47113
rect 64259 47085 64287 47113
rect 64321 47085 64349 47113
rect 64383 47085 64411 47113
rect 64197 47023 64225 47051
rect 64259 47023 64287 47051
rect 64321 47023 64349 47051
rect 64383 47023 64411 47051
rect 64197 46961 64225 46989
rect 64259 46961 64287 46989
rect 64321 46961 64349 46989
rect 64383 46961 64411 46989
rect 64197 38147 64225 38175
rect 64259 38147 64287 38175
rect 64321 38147 64349 38175
rect 64383 38147 64411 38175
rect 64197 38085 64225 38113
rect 64259 38085 64287 38113
rect 64321 38085 64349 38113
rect 64383 38085 64411 38113
rect 64197 38023 64225 38051
rect 64259 38023 64287 38051
rect 64321 38023 64349 38051
rect 64383 38023 64411 38051
rect 64197 37961 64225 37989
rect 64259 37961 64287 37989
rect 64321 37961 64349 37989
rect 64383 37961 64411 37989
rect 64197 29147 64225 29175
rect 64259 29147 64287 29175
rect 64321 29147 64349 29175
rect 64383 29147 64411 29175
rect 64197 29085 64225 29113
rect 64259 29085 64287 29113
rect 64321 29085 64349 29113
rect 64383 29085 64411 29113
rect 64197 29023 64225 29051
rect 64259 29023 64287 29051
rect 64321 29023 64349 29051
rect 64383 29023 64411 29051
rect 64197 28961 64225 28989
rect 64259 28961 64287 28989
rect 64321 28961 64349 28989
rect 64383 28961 64411 28989
rect 64197 20147 64225 20175
rect 64259 20147 64287 20175
rect 64321 20147 64349 20175
rect 64383 20147 64411 20175
rect 64197 20085 64225 20113
rect 64259 20085 64287 20113
rect 64321 20085 64349 20113
rect 64383 20085 64411 20113
rect 64197 20023 64225 20051
rect 64259 20023 64287 20051
rect 64321 20023 64349 20051
rect 64383 20023 64411 20051
rect 64197 19961 64225 19989
rect 64259 19961 64287 19989
rect 64321 19961 64349 19989
rect 64383 19961 64411 19989
rect 64197 11147 64225 11175
rect 64259 11147 64287 11175
rect 64321 11147 64349 11175
rect 64383 11147 64411 11175
rect 64197 11085 64225 11113
rect 64259 11085 64287 11113
rect 64321 11085 64349 11113
rect 64383 11085 64411 11113
rect 64197 11023 64225 11051
rect 64259 11023 64287 11051
rect 64321 11023 64349 11051
rect 64383 11023 64411 11051
rect 64197 10961 64225 10989
rect 64259 10961 64287 10989
rect 64321 10961 64349 10989
rect 64383 10961 64411 10989
rect 64197 2147 64225 2175
rect 64259 2147 64287 2175
rect 64321 2147 64349 2175
rect 64383 2147 64411 2175
rect 64197 2085 64225 2113
rect 64259 2085 64287 2113
rect 64321 2085 64349 2113
rect 64383 2085 64411 2113
rect 64197 2023 64225 2051
rect 64259 2023 64287 2051
rect 64321 2023 64349 2051
rect 64383 2023 64411 2051
rect 64197 1961 64225 1989
rect 64259 1961 64287 1989
rect 64321 1961 64349 1989
rect 64383 1961 64411 1989
rect 64197 -108 64225 -80
rect 64259 -108 64287 -80
rect 64321 -108 64349 -80
rect 64383 -108 64411 -80
rect 64197 -170 64225 -142
rect 64259 -170 64287 -142
rect 64321 -170 64349 -142
rect 64383 -170 64411 -142
rect 64197 -232 64225 -204
rect 64259 -232 64287 -204
rect 64321 -232 64349 -204
rect 64383 -232 64411 -204
rect 64197 -294 64225 -266
rect 64259 -294 64287 -266
rect 64321 -294 64349 -266
rect 64383 -294 64411 -266
rect 66057 68147 66085 68175
rect 66119 68147 66147 68175
rect 66181 68147 66209 68175
rect 66243 68147 66271 68175
rect 66057 68085 66085 68113
rect 66119 68085 66147 68113
rect 66181 68085 66209 68113
rect 66243 68085 66271 68113
rect 66057 68023 66085 68051
rect 66119 68023 66147 68051
rect 66181 68023 66209 68051
rect 66243 68023 66271 68051
rect 66057 67961 66085 67989
rect 66119 67961 66147 67989
rect 66181 67961 66209 67989
rect 66243 67961 66271 67989
rect 66057 59147 66085 59175
rect 66119 59147 66147 59175
rect 66181 59147 66209 59175
rect 66243 59147 66271 59175
rect 66057 59085 66085 59113
rect 66119 59085 66147 59113
rect 66181 59085 66209 59113
rect 66243 59085 66271 59113
rect 66057 59023 66085 59051
rect 66119 59023 66147 59051
rect 66181 59023 66209 59051
rect 66243 59023 66271 59051
rect 66057 58961 66085 58989
rect 66119 58961 66147 58989
rect 66181 58961 66209 58989
rect 66243 58961 66271 58989
rect 66057 50147 66085 50175
rect 66119 50147 66147 50175
rect 66181 50147 66209 50175
rect 66243 50147 66271 50175
rect 66057 50085 66085 50113
rect 66119 50085 66147 50113
rect 66181 50085 66209 50113
rect 66243 50085 66271 50113
rect 66057 50023 66085 50051
rect 66119 50023 66147 50051
rect 66181 50023 66209 50051
rect 66243 50023 66271 50051
rect 66057 49961 66085 49989
rect 66119 49961 66147 49989
rect 66181 49961 66209 49989
rect 66243 49961 66271 49989
rect 66057 41147 66085 41175
rect 66119 41147 66147 41175
rect 66181 41147 66209 41175
rect 66243 41147 66271 41175
rect 66057 41085 66085 41113
rect 66119 41085 66147 41113
rect 66181 41085 66209 41113
rect 66243 41085 66271 41113
rect 66057 41023 66085 41051
rect 66119 41023 66147 41051
rect 66181 41023 66209 41051
rect 66243 41023 66271 41051
rect 66057 40961 66085 40989
rect 66119 40961 66147 40989
rect 66181 40961 66209 40989
rect 66243 40961 66271 40989
rect 66057 32147 66085 32175
rect 66119 32147 66147 32175
rect 66181 32147 66209 32175
rect 66243 32147 66271 32175
rect 66057 32085 66085 32113
rect 66119 32085 66147 32113
rect 66181 32085 66209 32113
rect 66243 32085 66271 32113
rect 66057 32023 66085 32051
rect 66119 32023 66147 32051
rect 66181 32023 66209 32051
rect 66243 32023 66271 32051
rect 66057 31961 66085 31989
rect 66119 31961 66147 31989
rect 66181 31961 66209 31989
rect 66243 31961 66271 31989
rect 66057 23147 66085 23175
rect 66119 23147 66147 23175
rect 66181 23147 66209 23175
rect 66243 23147 66271 23175
rect 66057 23085 66085 23113
rect 66119 23085 66147 23113
rect 66181 23085 66209 23113
rect 66243 23085 66271 23113
rect 66057 23023 66085 23051
rect 66119 23023 66147 23051
rect 66181 23023 66209 23051
rect 66243 23023 66271 23051
rect 66057 22961 66085 22989
rect 66119 22961 66147 22989
rect 66181 22961 66209 22989
rect 66243 22961 66271 22989
rect 66057 14147 66085 14175
rect 66119 14147 66147 14175
rect 66181 14147 66209 14175
rect 66243 14147 66271 14175
rect 66057 14085 66085 14113
rect 66119 14085 66147 14113
rect 66181 14085 66209 14113
rect 66243 14085 66271 14113
rect 66057 14023 66085 14051
rect 66119 14023 66147 14051
rect 66181 14023 66209 14051
rect 66243 14023 66271 14051
rect 66057 13961 66085 13989
rect 66119 13961 66147 13989
rect 66181 13961 66209 13989
rect 66243 13961 66271 13989
rect 66057 5147 66085 5175
rect 66119 5147 66147 5175
rect 66181 5147 66209 5175
rect 66243 5147 66271 5175
rect 66057 5085 66085 5113
rect 66119 5085 66147 5113
rect 66181 5085 66209 5113
rect 66243 5085 66271 5113
rect 66057 5023 66085 5051
rect 66119 5023 66147 5051
rect 66181 5023 66209 5051
rect 66243 5023 66271 5051
rect 66057 4961 66085 4989
rect 66119 4961 66147 4989
rect 66181 4961 66209 4989
rect 66243 4961 66271 4989
rect 66057 -588 66085 -560
rect 66119 -588 66147 -560
rect 66181 -588 66209 -560
rect 66243 -588 66271 -560
rect 66057 -650 66085 -622
rect 66119 -650 66147 -622
rect 66181 -650 66209 -622
rect 66243 -650 66271 -622
rect 66057 -712 66085 -684
rect 66119 -712 66147 -684
rect 66181 -712 66209 -684
rect 66243 -712 66271 -684
rect 66057 -774 66085 -746
rect 66119 -774 66147 -746
rect 66181 -774 66209 -746
rect 66243 -774 66271 -746
rect 79557 74147 79585 74175
rect 79619 74147 79647 74175
rect 79681 74147 79709 74175
rect 79743 74147 79771 74175
rect 79557 74085 79585 74113
rect 79619 74085 79647 74113
rect 79681 74085 79709 74113
rect 79743 74085 79771 74113
rect 79557 74023 79585 74051
rect 79619 74023 79647 74051
rect 79681 74023 79709 74051
rect 79743 74023 79771 74051
rect 79557 73961 79585 73989
rect 79619 73961 79647 73989
rect 79681 73961 79709 73989
rect 79743 73961 79771 73989
rect 79557 65147 79585 65175
rect 79619 65147 79647 65175
rect 79681 65147 79709 65175
rect 79743 65147 79771 65175
rect 79557 65085 79585 65113
rect 79619 65085 79647 65113
rect 79681 65085 79709 65113
rect 79743 65085 79771 65113
rect 79557 65023 79585 65051
rect 79619 65023 79647 65051
rect 79681 65023 79709 65051
rect 79743 65023 79771 65051
rect 79557 64961 79585 64989
rect 79619 64961 79647 64989
rect 79681 64961 79709 64989
rect 79743 64961 79771 64989
rect 79557 56147 79585 56175
rect 79619 56147 79647 56175
rect 79681 56147 79709 56175
rect 79743 56147 79771 56175
rect 79557 56085 79585 56113
rect 79619 56085 79647 56113
rect 79681 56085 79709 56113
rect 79743 56085 79771 56113
rect 79557 56023 79585 56051
rect 79619 56023 79647 56051
rect 79681 56023 79709 56051
rect 79743 56023 79771 56051
rect 79557 55961 79585 55989
rect 79619 55961 79647 55989
rect 79681 55961 79709 55989
rect 79743 55961 79771 55989
rect 79557 47147 79585 47175
rect 79619 47147 79647 47175
rect 79681 47147 79709 47175
rect 79743 47147 79771 47175
rect 79557 47085 79585 47113
rect 79619 47085 79647 47113
rect 79681 47085 79709 47113
rect 79743 47085 79771 47113
rect 79557 47023 79585 47051
rect 79619 47023 79647 47051
rect 79681 47023 79709 47051
rect 79743 47023 79771 47051
rect 79557 46961 79585 46989
rect 79619 46961 79647 46989
rect 79681 46961 79709 46989
rect 79743 46961 79771 46989
rect 79557 38147 79585 38175
rect 79619 38147 79647 38175
rect 79681 38147 79709 38175
rect 79743 38147 79771 38175
rect 79557 38085 79585 38113
rect 79619 38085 79647 38113
rect 79681 38085 79709 38113
rect 79743 38085 79771 38113
rect 79557 38023 79585 38051
rect 79619 38023 79647 38051
rect 79681 38023 79709 38051
rect 79743 38023 79771 38051
rect 79557 37961 79585 37989
rect 79619 37961 79647 37989
rect 79681 37961 79709 37989
rect 79743 37961 79771 37989
rect 79557 29147 79585 29175
rect 79619 29147 79647 29175
rect 79681 29147 79709 29175
rect 79743 29147 79771 29175
rect 79557 29085 79585 29113
rect 79619 29085 79647 29113
rect 79681 29085 79709 29113
rect 79743 29085 79771 29113
rect 79557 29023 79585 29051
rect 79619 29023 79647 29051
rect 79681 29023 79709 29051
rect 79743 29023 79771 29051
rect 79557 28961 79585 28989
rect 79619 28961 79647 28989
rect 79681 28961 79709 28989
rect 79743 28961 79771 28989
rect 79557 20147 79585 20175
rect 79619 20147 79647 20175
rect 79681 20147 79709 20175
rect 79743 20147 79771 20175
rect 79557 20085 79585 20113
rect 79619 20085 79647 20113
rect 79681 20085 79709 20113
rect 79743 20085 79771 20113
rect 79557 20023 79585 20051
rect 79619 20023 79647 20051
rect 79681 20023 79709 20051
rect 79743 20023 79771 20051
rect 79557 19961 79585 19989
rect 79619 19961 79647 19989
rect 79681 19961 79709 19989
rect 79743 19961 79771 19989
rect 79557 11147 79585 11175
rect 79619 11147 79647 11175
rect 79681 11147 79709 11175
rect 79743 11147 79771 11175
rect 79557 11085 79585 11113
rect 79619 11085 79647 11113
rect 79681 11085 79709 11113
rect 79743 11085 79771 11113
rect 79557 11023 79585 11051
rect 79619 11023 79647 11051
rect 79681 11023 79709 11051
rect 79743 11023 79771 11051
rect 79557 10961 79585 10989
rect 79619 10961 79647 10989
rect 79681 10961 79709 10989
rect 79743 10961 79771 10989
rect 79557 2147 79585 2175
rect 79619 2147 79647 2175
rect 79681 2147 79709 2175
rect 79743 2147 79771 2175
rect 79557 2085 79585 2113
rect 79619 2085 79647 2113
rect 79681 2085 79709 2113
rect 79743 2085 79771 2113
rect 79557 2023 79585 2051
rect 79619 2023 79647 2051
rect 79681 2023 79709 2051
rect 79743 2023 79771 2051
rect 79557 1961 79585 1989
rect 79619 1961 79647 1989
rect 79681 1961 79709 1989
rect 79743 1961 79771 1989
rect 79557 -108 79585 -80
rect 79619 -108 79647 -80
rect 79681 -108 79709 -80
rect 79743 -108 79771 -80
rect 79557 -170 79585 -142
rect 79619 -170 79647 -142
rect 79681 -170 79709 -142
rect 79743 -170 79771 -142
rect 79557 -232 79585 -204
rect 79619 -232 79647 -204
rect 79681 -232 79709 -204
rect 79743 -232 79771 -204
rect 79557 -294 79585 -266
rect 79619 -294 79647 -266
rect 79681 -294 79709 -266
rect 79743 -294 79771 -266
rect 81417 167147 81445 167175
rect 81479 167147 81507 167175
rect 81541 167147 81569 167175
rect 81603 167147 81631 167175
rect 81417 167085 81445 167113
rect 81479 167085 81507 167113
rect 81541 167085 81569 167113
rect 81603 167085 81631 167113
rect 81417 167023 81445 167051
rect 81479 167023 81507 167051
rect 81541 167023 81569 167051
rect 81603 167023 81631 167051
rect 81417 166961 81445 166989
rect 81479 166961 81507 166989
rect 81541 166961 81569 166989
rect 81603 166961 81631 166989
rect 94917 164147 94945 164175
rect 94979 164147 95007 164175
rect 95041 164147 95069 164175
rect 95103 164147 95131 164175
rect 94917 164085 94945 164113
rect 94979 164085 95007 164113
rect 95041 164085 95069 164113
rect 95103 164085 95131 164113
rect 94917 164023 94945 164051
rect 94979 164023 95007 164051
rect 95041 164023 95069 164051
rect 95103 164023 95131 164051
rect 94917 163961 94945 163989
rect 94979 163961 95007 163989
rect 95041 163961 95069 163989
rect 95103 163961 95131 163989
rect 81417 158147 81445 158175
rect 81479 158147 81507 158175
rect 81541 158147 81569 158175
rect 81603 158147 81631 158175
rect 81417 158085 81445 158113
rect 81479 158085 81507 158113
rect 81541 158085 81569 158113
rect 81603 158085 81631 158113
rect 81417 158023 81445 158051
rect 81479 158023 81507 158051
rect 81541 158023 81569 158051
rect 81603 158023 81631 158051
rect 81417 157961 81445 157989
rect 81479 157961 81507 157989
rect 81541 157961 81569 157989
rect 81603 157961 81631 157989
rect 86019 158147 86047 158175
rect 86081 158147 86109 158175
rect 86019 158085 86047 158113
rect 86081 158085 86109 158113
rect 86019 158023 86047 158051
rect 86081 158023 86109 158051
rect 86019 157961 86047 157989
rect 86081 157961 86109 157989
rect 93699 155147 93727 155175
rect 93761 155147 93789 155175
rect 93699 155085 93727 155113
rect 93761 155085 93789 155113
rect 93699 155023 93727 155051
rect 93761 155023 93789 155051
rect 93699 154961 93727 154989
rect 93761 154961 93789 154989
rect 94917 155147 94945 155175
rect 94979 155147 95007 155175
rect 95041 155147 95069 155175
rect 95103 155147 95131 155175
rect 94917 155085 94945 155113
rect 94979 155085 95007 155113
rect 95041 155085 95069 155113
rect 95103 155085 95131 155113
rect 94917 155023 94945 155051
rect 94979 155023 95007 155051
rect 95041 155023 95069 155051
rect 95103 155023 95131 155051
rect 94917 154961 94945 154989
rect 94979 154961 95007 154989
rect 95041 154961 95069 154989
rect 95103 154961 95131 154989
rect 81417 149147 81445 149175
rect 81479 149147 81507 149175
rect 81541 149147 81569 149175
rect 81603 149147 81631 149175
rect 81417 149085 81445 149113
rect 81479 149085 81507 149113
rect 81541 149085 81569 149113
rect 81603 149085 81631 149113
rect 81417 149023 81445 149051
rect 81479 149023 81507 149051
rect 81541 149023 81569 149051
rect 81603 149023 81631 149051
rect 81417 148961 81445 148989
rect 81479 148961 81507 148989
rect 81541 148961 81569 148989
rect 81603 148961 81631 148989
rect 86019 149147 86047 149175
rect 86081 149147 86109 149175
rect 86019 149085 86047 149113
rect 86081 149085 86109 149113
rect 86019 149023 86047 149051
rect 86081 149023 86109 149051
rect 86019 148961 86047 148989
rect 86081 148961 86109 148989
rect 93699 146147 93727 146175
rect 93761 146147 93789 146175
rect 93699 146085 93727 146113
rect 93761 146085 93789 146113
rect 93699 146023 93727 146051
rect 93761 146023 93789 146051
rect 93699 145961 93727 145989
rect 93761 145961 93789 145989
rect 94917 146147 94945 146175
rect 94979 146147 95007 146175
rect 95041 146147 95069 146175
rect 95103 146147 95131 146175
rect 94917 146085 94945 146113
rect 94979 146085 95007 146113
rect 95041 146085 95069 146113
rect 95103 146085 95131 146113
rect 94917 146023 94945 146051
rect 94979 146023 95007 146051
rect 95041 146023 95069 146051
rect 95103 146023 95131 146051
rect 94917 145961 94945 145989
rect 94979 145961 95007 145989
rect 95041 145961 95069 145989
rect 95103 145961 95131 145989
rect 81417 140147 81445 140175
rect 81479 140147 81507 140175
rect 81541 140147 81569 140175
rect 81603 140147 81631 140175
rect 81417 140085 81445 140113
rect 81479 140085 81507 140113
rect 81541 140085 81569 140113
rect 81603 140085 81631 140113
rect 81417 140023 81445 140051
rect 81479 140023 81507 140051
rect 81541 140023 81569 140051
rect 81603 140023 81631 140051
rect 81417 139961 81445 139989
rect 81479 139961 81507 139989
rect 81541 139961 81569 139989
rect 81603 139961 81631 139989
rect 86019 140147 86047 140175
rect 86081 140147 86109 140175
rect 86019 140085 86047 140113
rect 86081 140085 86109 140113
rect 86019 140023 86047 140051
rect 86081 140023 86109 140051
rect 86019 139961 86047 139989
rect 86081 139961 86109 139989
rect 93699 137147 93727 137175
rect 93761 137147 93789 137175
rect 93699 137085 93727 137113
rect 93761 137085 93789 137113
rect 93699 137023 93727 137051
rect 93761 137023 93789 137051
rect 93699 136961 93727 136989
rect 93761 136961 93789 136989
rect 94917 137147 94945 137175
rect 94979 137147 95007 137175
rect 95041 137147 95069 137175
rect 95103 137147 95131 137175
rect 94917 137085 94945 137113
rect 94979 137085 95007 137113
rect 95041 137085 95069 137113
rect 95103 137085 95131 137113
rect 94917 137023 94945 137051
rect 94979 137023 95007 137051
rect 95041 137023 95069 137051
rect 95103 137023 95131 137051
rect 94917 136961 94945 136989
rect 94979 136961 95007 136989
rect 95041 136961 95069 136989
rect 95103 136961 95131 136989
rect 81417 131147 81445 131175
rect 81479 131147 81507 131175
rect 81541 131147 81569 131175
rect 81603 131147 81631 131175
rect 81417 131085 81445 131113
rect 81479 131085 81507 131113
rect 81541 131085 81569 131113
rect 81603 131085 81631 131113
rect 81417 131023 81445 131051
rect 81479 131023 81507 131051
rect 81541 131023 81569 131051
rect 81603 131023 81631 131051
rect 81417 130961 81445 130989
rect 81479 130961 81507 130989
rect 81541 130961 81569 130989
rect 81603 130961 81631 130989
rect 81417 122147 81445 122175
rect 81479 122147 81507 122175
rect 81541 122147 81569 122175
rect 81603 122147 81631 122175
rect 81417 122085 81445 122113
rect 81479 122085 81507 122113
rect 81541 122085 81569 122113
rect 81603 122085 81631 122113
rect 81417 122023 81445 122051
rect 81479 122023 81507 122051
rect 81541 122023 81569 122051
rect 81603 122023 81631 122051
rect 81417 121961 81445 121989
rect 81479 121961 81507 121989
rect 81541 121961 81569 121989
rect 81603 121961 81631 121989
rect 81417 113147 81445 113175
rect 81479 113147 81507 113175
rect 81541 113147 81569 113175
rect 81603 113147 81631 113175
rect 81417 113085 81445 113113
rect 81479 113085 81507 113113
rect 81541 113085 81569 113113
rect 81603 113085 81631 113113
rect 81417 113023 81445 113051
rect 81479 113023 81507 113051
rect 81541 113023 81569 113051
rect 81603 113023 81631 113051
rect 81417 112961 81445 112989
rect 81479 112961 81507 112989
rect 81541 112961 81569 112989
rect 81603 112961 81631 112989
rect 81417 104147 81445 104175
rect 81479 104147 81507 104175
rect 81541 104147 81569 104175
rect 81603 104147 81631 104175
rect 81417 104085 81445 104113
rect 81479 104085 81507 104113
rect 81541 104085 81569 104113
rect 81603 104085 81631 104113
rect 81417 104023 81445 104051
rect 81479 104023 81507 104051
rect 81541 104023 81569 104051
rect 81603 104023 81631 104051
rect 81417 103961 81445 103989
rect 81479 103961 81507 103989
rect 81541 103961 81569 103989
rect 81603 103961 81631 103989
rect 94917 128147 94945 128175
rect 94979 128147 95007 128175
rect 95041 128147 95069 128175
rect 95103 128147 95131 128175
rect 94917 128085 94945 128113
rect 94979 128085 95007 128113
rect 95041 128085 95069 128113
rect 95103 128085 95131 128113
rect 94917 128023 94945 128051
rect 94979 128023 95007 128051
rect 95041 128023 95069 128051
rect 95103 128023 95131 128051
rect 94917 127961 94945 127989
rect 94979 127961 95007 127989
rect 95041 127961 95069 127989
rect 95103 127961 95131 127989
rect 94917 119147 94945 119175
rect 94979 119147 95007 119175
rect 95041 119147 95069 119175
rect 95103 119147 95131 119175
rect 94917 119085 94945 119113
rect 94979 119085 95007 119113
rect 95041 119085 95069 119113
rect 95103 119085 95131 119113
rect 94917 119023 94945 119051
rect 94979 119023 95007 119051
rect 95041 119023 95069 119051
rect 95103 119023 95131 119051
rect 94917 118961 94945 118989
rect 94979 118961 95007 118989
rect 95041 118961 95069 118989
rect 95103 118961 95131 118989
rect 94917 110147 94945 110175
rect 94979 110147 95007 110175
rect 95041 110147 95069 110175
rect 95103 110147 95131 110175
rect 94917 110085 94945 110113
rect 94979 110085 95007 110113
rect 95041 110085 95069 110113
rect 95103 110085 95131 110113
rect 94917 110023 94945 110051
rect 94979 110023 95007 110051
rect 95041 110023 95069 110051
rect 95103 110023 95131 110051
rect 94917 109961 94945 109989
rect 94979 109961 95007 109989
rect 95041 109961 95069 109989
rect 95103 109961 95131 109989
rect 93059 101147 93087 101175
rect 93121 101147 93149 101175
rect 93059 101085 93087 101113
rect 93121 101085 93149 101113
rect 93059 101023 93087 101051
rect 93121 101023 93149 101051
rect 93059 100961 93087 100989
rect 93121 100961 93149 100989
rect 94917 101147 94945 101175
rect 94979 101147 95007 101175
rect 95041 101147 95069 101175
rect 95103 101147 95131 101175
rect 94917 101085 94945 101113
rect 94979 101085 95007 101113
rect 95041 101085 95069 101113
rect 95103 101085 95131 101113
rect 94917 101023 94945 101051
rect 94979 101023 95007 101051
rect 95041 101023 95069 101051
rect 95103 101023 95131 101051
rect 94917 100961 94945 100989
rect 94979 100961 95007 100989
rect 95041 100961 95069 100989
rect 95103 100961 95131 100989
rect 81417 95147 81445 95175
rect 81479 95147 81507 95175
rect 81541 95147 81569 95175
rect 81603 95147 81631 95175
rect 81417 95085 81445 95113
rect 81479 95085 81507 95113
rect 81541 95085 81569 95113
rect 81603 95085 81631 95113
rect 81417 95023 81445 95051
rect 81479 95023 81507 95051
rect 81541 95023 81569 95051
rect 81603 95023 81631 95051
rect 81417 94961 81445 94989
rect 81479 94961 81507 94989
rect 81541 94961 81569 94989
rect 81603 94961 81631 94989
rect 85379 95147 85407 95175
rect 85441 95147 85469 95175
rect 85379 95085 85407 95113
rect 85441 95085 85469 95113
rect 85379 95023 85407 95051
rect 85441 95023 85469 95051
rect 85379 94961 85407 94989
rect 85441 94961 85469 94989
rect 93059 92147 93087 92175
rect 93121 92147 93149 92175
rect 93059 92085 93087 92113
rect 93121 92085 93149 92113
rect 93059 92023 93087 92051
rect 93121 92023 93149 92051
rect 93059 91961 93087 91989
rect 93121 91961 93149 91989
rect 94917 92147 94945 92175
rect 94979 92147 95007 92175
rect 95041 92147 95069 92175
rect 95103 92147 95131 92175
rect 94917 92085 94945 92113
rect 94979 92085 95007 92113
rect 95041 92085 95069 92113
rect 95103 92085 95131 92113
rect 94917 92023 94945 92051
rect 94979 92023 95007 92051
rect 95041 92023 95069 92051
rect 95103 92023 95131 92051
rect 94917 91961 94945 91989
rect 94979 91961 95007 91989
rect 95041 91961 95069 91989
rect 95103 91961 95131 91989
rect 81417 86147 81445 86175
rect 81479 86147 81507 86175
rect 81541 86147 81569 86175
rect 81603 86147 81631 86175
rect 81417 86085 81445 86113
rect 81479 86085 81507 86113
rect 81541 86085 81569 86113
rect 81603 86085 81631 86113
rect 81417 86023 81445 86051
rect 81479 86023 81507 86051
rect 81541 86023 81569 86051
rect 81603 86023 81631 86051
rect 81417 85961 81445 85989
rect 81479 85961 81507 85989
rect 81541 85961 81569 85989
rect 81603 85961 81631 85989
rect 85379 86147 85407 86175
rect 85441 86147 85469 86175
rect 85379 86085 85407 86113
rect 85441 86085 85469 86113
rect 85379 86023 85407 86051
rect 85441 86023 85469 86051
rect 85379 85961 85407 85989
rect 85441 85961 85469 85989
rect 93059 83147 93087 83175
rect 93121 83147 93149 83175
rect 93059 83085 93087 83113
rect 93121 83085 93149 83113
rect 93059 83023 93087 83051
rect 93121 83023 93149 83051
rect 93059 82961 93087 82989
rect 93121 82961 93149 82989
rect 94917 83147 94945 83175
rect 94979 83147 95007 83175
rect 95041 83147 95069 83175
rect 95103 83147 95131 83175
rect 94917 83085 94945 83113
rect 94979 83085 95007 83113
rect 95041 83085 95069 83113
rect 95103 83085 95131 83113
rect 94917 83023 94945 83051
rect 94979 83023 95007 83051
rect 95041 83023 95069 83051
rect 95103 83023 95131 83051
rect 94917 82961 94945 82989
rect 94979 82961 95007 82989
rect 95041 82961 95069 82989
rect 95103 82961 95131 82989
rect 81417 77147 81445 77175
rect 81479 77147 81507 77175
rect 81541 77147 81569 77175
rect 81603 77147 81631 77175
rect 81417 77085 81445 77113
rect 81479 77085 81507 77113
rect 81541 77085 81569 77113
rect 81603 77085 81631 77113
rect 81417 77023 81445 77051
rect 81479 77023 81507 77051
rect 81541 77023 81569 77051
rect 81603 77023 81631 77051
rect 81417 76961 81445 76989
rect 81479 76961 81507 76989
rect 81541 76961 81569 76989
rect 81603 76961 81631 76989
rect 85379 77147 85407 77175
rect 85441 77147 85469 77175
rect 85379 77085 85407 77113
rect 85441 77085 85469 77113
rect 85379 77023 85407 77051
rect 85441 77023 85469 77051
rect 85379 76961 85407 76989
rect 85441 76961 85469 76989
rect 81417 68147 81445 68175
rect 81479 68147 81507 68175
rect 81541 68147 81569 68175
rect 81603 68147 81631 68175
rect 81417 68085 81445 68113
rect 81479 68085 81507 68113
rect 81541 68085 81569 68113
rect 81603 68085 81631 68113
rect 81417 68023 81445 68051
rect 81479 68023 81507 68051
rect 81541 68023 81569 68051
rect 81603 68023 81631 68051
rect 81417 67961 81445 67989
rect 81479 67961 81507 67989
rect 81541 67961 81569 67989
rect 81603 67961 81631 67989
rect 81417 59147 81445 59175
rect 81479 59147 81507 59175
rect 81541 59147 81569 59175
rect 81603 59147 81631 59175
rect 81417 59085 81445 59113
rect 81479 59085 81507 59113
rect 81541 59085 81569 59113
rect 81603 59085 81631 59113
rect 81417 59023 81445 59051
rect 81479 59023 81507 59051
rect 81541 59023 81569 59051
rect 81603 59023 81631 59051
rect 81417 58961 81445 58989
rect 81479 58961 81507 58989
rect 81541 58961 81569 58989
rect 81603 58961 81631 58989
rect 81417 50147 81445 50175
rect 81479 50147 81507 50175
rect 81541 50147 81569 50175
rect 81603 50147 81631 50175
rect 81417 50085 81445 50113
rect 81479 50085 81507 50113
rect 81541 50085 81569 50113
rect 81603 50085 81631 50113
rect 81417 50023 81445 50051
rect 81479 50023 81507 50051
rect 81541 50023 81569 50051
rect 81603 50023 81631 50051
rect 81417 49961 81445 49989
rect 81479 49961 81507 49989
rect 81541 49961 81569 49989
rect 81603 49961 81631 49989
rect 81417 41147 81445 41175
rect 81479 41147 81507 41175
rect 81541 41147 81569 41175
rect 81603 41147 81631 41175
rect 81417 41085 81445 41113
rect 81479 41085 81507 41113
rect 81541 41085 81569 41113
rect 81603 41085 81631 41113
rect 81417 41023 81445 41051
rect 81479 41023 81507 41051
rect 81541 41023 81569 41051
rect 81603 41023 81631 41051
rect 81417 40961 81445 40989
rect 81479 40961 81507 40989
rect 81541 40961 81569 40989
rect 81603 40961 81631 40989
rect 81417 32147 81445 32175
rect 81479 32147 81507 32175
rect 81541 32147 81569 32175
rect 81603 32147 81631 32175
rect 81417 32085 81445 32113
rect 81479 32085 81507 32113
rect 81541 32085 81569 32113
rect 81603 32085 81631 32113
rect 81417 32023 81445 32051
rect 81479 32023 81507 32051
rect 81541 32023 81569 32051
rect 81603 32023 81631 32051
rect 81417 31961 81445 31989
rect 81479 31961 81507 31989
rect 81541 31961 81569 31989
rect 81603 31961 81631 31989
rect 81417 23147 81445 23175
rect 81479 23147 81507 23175
rect 81541 23147 81569 23175
rect 81603 23147 81631 23175
rect 81417 23085 81445 23113
rect 81479 23085 81507 23113
rect 81541 23085 81569 23113
rect 81603 23085 81631 23113
rect 81417 23023 81445 23051
rect 81479 23023 81507 23051
rect 81541 23023 81569 23051
rect 81603 23023 81631 23051
rect 81417 22961 81445 22989
rect 81479 22961 81507 22989
rect 81541 22961 81569 22989
rect 81603 22961 81631 22989
rect 81417 14147 81445 14175
rect 81479 14147 81507 14175
rect 81541 14147 81569 14175
rect 81603 14147 81631 14175
rect 81417 14085 81445 14113
rect 81479 14085 81507 14113
rect 81541 14085 81569 14113
rect 81603 14085 81631 14113
rect 81417 14023 81445 14051
rect 81479 14023 81507 14051
rect 81541 14023 81569 14051
rect 81603 14023 81631 14051
rect 81417 13961 81445 13989
rect 81479 13961 81507 13989
rect 81541 13961 81569 13989
rect 81603 13961 81631 13989
rect 81417 5147 81445 5175
rect 81479 5147 81507 5175
rect 81541 5147 81569 5175
rect 81603 5147 81631 5175
rect 81417 5085 81445 5113
rect 81479 5085 81507 5113
rect 81541 5085 81569 5113
rect 81603 5085 81631 5113
rect 81417 5023 81445 5051
rect 81479 5023 81507 5051
rect 81541 5023 81569 5051
rect 81603 5023 81631 5051
rect 81417 4961 81445 4989
rect 81479 4961 81507 4989
rect 81541 4961 81569 4989
rect 81603 4961 81631 4989
rect 81417 -588 81445 -560
rect 81479 -588 81507 -560
rect 81541 -588 81569 -560
rect 81603 -588 81631 -560
rect 81417 -650 81445 -622
rect 81479 -650 81507 -622
rect 81541 -650 81569 -622
rect 81603 -650 81631 -622
rect 81417 -712 81445 -684
rect 81479 -712 81507 -684
rect 81541 -712 81569 -684
rect 81603 -712 81631 -684
rect 81417 -774 81445 -746
rect 81479 -774 81507 -746
rect 81541 -774 81569 -746
rect 81603 -774 81631 -746
rect 94917 74147 94945 74175
rect 94979 74147 95007 74175
rect 95041 74147 95069 74175
rect 95103 74147 95131 74175
rect 94917 74085 94945 74113
rect 94979 74085 95007 74113
rect 95041 74085 95069 74113
rect 95103 74085 95131 74113
rect 94917 74023 94945 74051
rect 94979 74023 95007 74051
rect 95041 74023 95069 74051
rect 95103 74023 95131 74051
rect 94917 73961 94945 73989
rect 94979 73961 95007 73989
rect 95041 73961 95069 73989
rect 95103 73961 95131 73989
rect 94917 65147 94945 65175
rect 94979 65147 95007 65175
rect 95041 65147 95069 65175
rect 95103 65147 95131 65175
rect 94917 65085 94945 65113
rect 94979 65085 95007 65113
rect 95041 65085 95069 65113
rect 95103 65085 95131 65113
rect 94917 65023 94945 65051
rect 94979 65023 95007 65051
rect 95041 65023 95069 65051
rect 95103 65023 95131 65051
rect 94917 64961 94945 64989
rect 94979 64961 95007 64989
rect 95041 64961 95069 64989
rect 95103 64961 95131 64989
rect 94917 56147 94945 56175
rect 94979 56147 95007 56175
rect 95041 56147 95069 56175
rect 95103 56147 95131 56175
rect 94917 56085 94945 56113
rect 94979 56085 95007 56113
rect 95041 56085 95069 56113
rect 95103 56085 95131 56113
rect 94917 56023 94945 56051
rect 94979 56023 95007 56051
rect 95041 56023 95069 56051
rect 95103 56023 95131 56051
rect 94917 55961 94945 55989
rect 94979 55961 95007 55989
rect 95041 55961 95069 55989
rect 95103 55961 95131 55989
rect 94917 47147 94945 47175
rect 94979 47147 95007 47175
rect 95041 47147 95069 47175
rect 95103 47147 95131 47175
rect 94917 47085 94945 47113
rect 94979 47085 95007 47113
rect 95041 47085 95069 47113
rect 95103 47085 95131 47113
rect 94917 47023 94945 47051
rect 94979 47023 95007 47051
rect 95041 47023 95069 47051
rect 95103 47023 95131 47051
rect 94917 46961 94945 46989
rect 94979 46961 95007 46989
rect 95041 46961 95069 46989
rect 95103 46961 95131 46989
rect 94917 38147 94945 38175
rect 94979 38147 95007 38175
rect 95041 38147 95069 38175
rect 95103 38147 95131 38175
rect 94917 38085 94945 38113
rect 94979 38085 95007 38113
rect 95041 38085 95069 38113
rect 95103 38085 95131 38113
rect 94917 38023 94945 38051
rect 94979 38023 95007 38051
rect 95041 38023 95069 38051
rect 95103 38023 95131 38051
rect 94917 37961 94945 37989
rect 94979 37961 95007 37989
rect 95041 37961 95069 37989
rect 95103 37961 95131 37989
rect 94917 29147 94945 29175
rect 94979 29147 95007 29175
rect 95041 29147 95069 29175
rect 95103 29147 95131 29175
rect 94917 29085 94945 29113
rect 94979 29085 95007 29113
rect 95041 29085 95069 29113
rect 95103 29085 95131 29113
rect 94917 29023 94945 29051
rect 94979 29023 95007 29051
rect 95041 29023 95069 29051
rect 95103 29023 95131 29051
rect 94917 28961 94945 28989
rect 94979 28961 95007 28989
rect 95041 28961 95069 28989
rect 95103 28961 95131 28989
rect 94917 20147 94945 20175
rect 94979 20147 95007 20175
rect 95041 20147 95069 20175
rect 95103 20147 95131 20175
rect 94917 20085 94945 20113
rect 94979 20085 95007 20113
rect 95041 20085 95069 20113
rect 95103 20085 95131 20113
rect 94917 20023 94945 20051
rect 94979 20023 95007 20051
rect 95041 20023 95069 20051
rect 95103 20023 95131 20051
rect 94917 19961 94945 19989
rect 94979 19961 95007 19989
rect 95041 19961 95069 19989
rect 95103 19961 95131 19989
rect 94917 11147 94945 11175
rect 94979 11147 95007 11175
rect 95041 11147 95069 11175
rect 95103 11147 95131 11175
rect 94917 11085 94945 11113
rect 94979 11085 95007 11113
rect 95041 11085 95069 11113
rect 95103 11085 95131 11113
rect 94917 11023 94945 11051
rect 94979 11023 95007 11051
rect 95041 11023 95069 11051
rect 95103 11023 95131 11051
rect 94917 10961 94945 10989
rect 94979 10961 95007 10989
rect 95041 10961 95069 10989
rect 95103 10961 95131 10989
rect 94917 2147 94945 2175
rect 94979 2147 95007 2175
rect 95041 2147 95069 2175
rect 95103 2147 95131 2175
rect 94917 2085 94945 2113
rect 94979 2085 95007 2113
rect 95041 2085 95069 2113
rect 95103 2085 95131 2113
rect 94917 2023 94945 2051
rect 94979 2023 95007 2051
rect 95041 2023 95069 2051
rect 95103 2023 95131 2051
rect 94917 1961 94945 1989
rect 94979 1961 95007 1989
rect 95041 1961 95069 1989
rect 95103 1961 95131 1989
rect 94917 -108 94945 -80
rect 94979 -108 95007 -80
rect 95041 -108 95069 -80
rect 95103 -108 95131 -80
rect 94917 -170 94945 -142
rect 94979 -170 95007 -142
rect 95041 -170 95069 -142
rect 95103 -170 95131 -142
rect 94917 -232 94945 -204
rect 94979 -232 95007 -204
rect 95041 -232 95069 -204
rect 95103 -232 95131 -204
rect 94917 -294 94945 -266
rect 94979 -294 95007 -266
rect 95041 -294 95069 -266
rect 95103 -294 95131 -266
rect 96777 299058 96805 299086
rect 96839 299058 96867 299086
rect 96901 299058 96929 299086
rect 96963 299058 96991 299086
rect 96777 298996 96805 299024
rect 96839 298996 96867 299024
rect 96901 298996 96929 299024
rect 96963 298996 96991 299024
rect 96777 298934 96805 298962
rect 96839 298934 96867 298962
rect 96901 298934 96929 298962
rect 96963 298934 96991 298962
rect 96777 298872 96805 298900
rect 96839 298872 96867 298900
rect 96901 298872 96929 298900
rect 96963 298872 96991 298900
rect 96777 293147 96805 293175
rect 96839 293147 96867 293175
rect 96901 293147 96929 293175
rect 96963 293147 96991 293175
rect 96777 293085 96805 293113
rect 96839 293085 96867 293113
rect 96901 293085 96929 293113
rect 96963 293085 96991 293113
rect 96777 293023 96805 293051
rect 96839 293023 96867 293051
rect 96901 293023 96929 293051
rect 96963 293023 96991 293051
rect 96777 292961 96805 292989
rect 96839 292961 96867 292989
rect 96901 292961 96929 292989
rect 96963 292961 96991 292989
rect 96777 284147 96805 284175
rect 96839 284147 96867 284175
rect 96901 284147 96929 284175
rect 96963 284147 96991 284175
rect 96777 284085 96805 284113
rect 96839 284085 96867 284113
rect 96901 284085 96929 284113
rect 96963 284085 96991 284113
rect 96777 284023 96805 284051
rect 96839 284023 96867 284051
rect 96901 284023 96929 284051
rect 96963 284023 96991 284051
rect 96777 283961 96805 283989
rect 96839 283961 96867 283989
rect 96901 283961 96929 283989
rect 96963 283961 96991 283989
rect 96777 275147 96805 275175
rect 96839 275147 96867 275175
rect 96901 275147 96929 275175
rect 96963 275147 96991 275175
rect 96777 275085 96805 275113
rect 96839 275085 96867 275113
rect 96901 275085 96929 275113
rect 96963 275085 96991 275113
rect 96777 275023 96805 275051
rect 96839 275023 96867 275051
rect 96901 275023 96929 275051
rect 96963 275023 96991 275051
rect 96777 274961 96805 274989
rect 96839 274961 96867 274989
rect 96901 274961 96929 274989
rect 96963 274961 96991 274989
rect 110277 298578 110305 298606
rect 110339 298578 110367 298606
rect 110401 298578 110429 298606
rect 110463 298578 110491 298606
rect 110277 298516 110305 298544
rect 110339 298516 110367 298544
rect 110401 298516 110429 298544
rect 110463 298516 110491 298544
rect 110277 298454 110305 298482
rect 110339 298454 110367 298482
rect 110401 298454 110429 298482
rect 110463 298454 110491 298482
rect 110277 298392 110305 298420
rect 110339 298392 110367 298420
rect 110401 298392 110429 298420
rect 110463 298392 110491 298420
rect 110277 290147 110305 290175
rect 110339 290147 110367 290175
rect 110401 290147 110429 290175
rect 110463 290147 110491 290175
rect 110277 290085 110305 290113
rect 110339 290085 110367 290113
rect 110401 290085 110429 290113
rect 110463 290085 110491 290113
rect 110277 290023 110305 290051
rect 110339 290023 110367 290051
rect 110401 290023 110429 290051
rect 110463 290023 110491 290051
rect 110277 289961 110305 289989
rect 110339 289961 110367 289989
rect 110401 289961 110429 289989
rect 110463 289961 110491 289989
rect 110277 281147 110305 281175
rect 110339 281147 110367 281175
rect 110401 281147 110429 281175
rect 110463 281147 110491 281175
rect 110277 281085 110305 281113
rect 110339 281085 110367 281113
rect 110401 281085 110429 281113
rect 110463 281085 110491 281113
rect 110277 281023 110305 281051
rect 110339 281023 110367 281051
rect 110401 281023 110429 281051
rect 110463 281023 110491 281051
rect 110277 280961 110305 280989
rect 110339 280961 110367 280989
rect 110401 280961 110429 280989
rect 110463 280961 110491 280989
rect 110277 272147 110305 272175
rect 110339 272147 110367 272175
rect 110401 272147 110429 272175
rect 110463 272147 110491 272175
rect 110277 272085 110305 272113
rect 110339 272085 110367 272113
rect 110401 272085 110429 272113
rect 110463 272085 110491 272113
rect 110277 272023 110305 272051
rect 110339 272023 110367 272051
rect 110401 272023 110429 272051
rect 110463 272023 110491 272051
rect 110277 271961 110305 271989
rect 110339 271961 110367 271989
rect 110401 271961 110429 271989
rect 110463 271961 110491 271989
rect 112137 299058 112165 299086
rect 112199 299058 112227 299086
rect 112261 299058 112289 299086
rect 112323 299058 112351 299086
rect 112137 298996 112165 299024
rect 112199 298996 112227 299024
rect 112261 298996 112289 299024
rect 112323 298996 112351 299024
rect 112137 298934 112165 298962
rect 112199 298934 112227 298962
rect 112261 298934 112289 298962
rect 112323 298934 112351 298962
rect 112137 298872 112165 298900
rect 112199 298872 112227 298900
rect 112261 298872 112289 298900
rect 112323 298872 112351 298900
rect 112137 293147 112165 293175
rect 112199 293147 112227 293175
rect 112261 293147 112289 293175
rect 112323 293147 112351 293175
rect 112137 293085 112165 293113
rect 112199 293085 112227 293113
rect 112261 293085 112289 293113
rect 112323 293085 112351 293113
rect 112137 293023 112165 293051
rect 112199 293023 112227 293051
rect 112261 293023 112289 293051
rect 112323 293023 112351 293051
rect 112137 292961 112165 292989
rect 112199 292961 112227 292989
rect 112261 292961 112289 292989
rect 112323 292961 112351 292989
rect 112137 284147 112165 284175
rect 112199 284147 112227 284175
rect 112261 284147 112289 284175
rect 112323 284147 112351 284175
rect 112137 284085 112165 284113
rect 112199 284085 112227 284113
rect 112261 284085 112289 284113
rect 112323 284085 112351 284113
rect 112137 284023 112165 284051
rect 112199 284023 112227 284051
rect 112261 284023 112289 284051
rect 112323 284023 112351 284051
rect 112137 283961 112165 283989
rect 112199 283961 112227 283989
rect 112261 283961 112289 283989
rect 112323 283961 112351 283989
rect 112137 275147 112165 275175
rect 112199 275147 112227 275175
rect 112261 275147 112289 275175
rect 112323 275147 112351 275175
rect 112137 275085 112165 275113
rect 112199 275085 112227 275113
rect 112261 275085 112289 275113
rect 112323 275085 112351 275113
rect 112137 275023 112165 275051
rect 112199 275023 112227 275051
rect 112261 275023 112289 275051
rect 112323 275023 112351 275051
rect 112137 274961 112165 274989
rect 112199 274961 112227 274989
rect 112261 274961 112289 274989
rect 112323 274961 112351 274989
rect 125637 298578 125665 298606
rect 125699 298578 125727 298606
rect 125761 298578 125789 298606
rect 125823 298578 125851 298606
rect 125637 298516 125665 298544
rect 125699 298516 125727 298544
rect 125761 298516 125789 298544
rect 125823 298516 125851 298544
rect 125637 298454 125665 298482
rect 125699 298454 125727 298482
rect 125761 298454 125789 298482
rect 125823 298454 125851 298482
rect 125637 298392 125665 298420
rect 125699 298392 125727 298420
rect 125761 298392 125789 298420
rect 125823 298392 125851 298420
rect 125637 290147 125665 290175
rect 125699 290147 125727 290175
rect 125761 290147 125789 290175
rect 125823 290147 125851 290175
rect 125637 290085 125665 290113
rect 125699 290085 125727 290113
rect 125761 290085 125789 290113
rect 125823 290085 125851 290113
rect 125637 290023 125665 290051
rect 125699 290023 125727 290051
rect 125761 290023 125789 290051
rect 125823 290023 125851 290051
rect 125637 289961 125665 289989
rect 125699 289961 125727 289989
rect 125761 289961 125789 289989
rect 125823 289961 125851 289989
rect 125637 281147 125665 281175
rect 125699 281147 125727 281175
rect 125761 281147 125789 281175
rect 125823 281147 125851 281175
rect 125637 281085 125665 281113
rect 125699 281085 125727 281113
rect 125761 281085 125789 281113
rect 125823 281085 125851 281113
rect 125637 281023 125665 281051
rect 125699 281023 125727 281051
rect 125761 281023 125789 281051
rect 125823 281023 125851 281051
rect 125637 280961 125665 280989
rect 125699 280961 125727 280989
rect 125761 280961 125789 280989
rect 125823 280961 125851 280989
rect 125637 272147 125665 272175
rect 125699 272147 125727 272175
rect 125761 272147 125789 272175
rect 125823 272147 125851 272175
rect 125637 272085 125665 272113
rect 125699 272085 125727 272113
rect 125761 272085 125789 272113
rect 125823 272085 125851 272113
rect 125637 272023 125665 272051
rect 125699 272023 125727 272051
rect 125761 272023 125789 272051
rect 125823 272023 125851 272051
rect 125637 271961 125665 271989
rect 125699 271961 125727 271989
rect 125761 271961 125789 271989
rect 125823 271961 125851 271989
rect 127497 299058 127525 299086
rect 127559 299058 127587 299086
rect 127621 299058 127649 299086
rect 127683 299058 127711 299086
rect 127497 298996 127525 299024
rect 127559 298996 127587 299024
rect 127621 298996 127649 299024
rect 127683 298996 127711 299024
rect 127497 298934 127525 298962
rect 127559 298934 127587 298962
rect 127621 298934 127649 298962
rect 127683 298934 127711 298962
rect 127497 298872 127525 298900
rect 127559 298872 127587 298900
rect 127621 298872 127649 298900
rect 127683 298872 127711 298900
rect 127497 293147 127525 293175
rect 127559 293147 127587 293175
rect 127621 293147 127649 293175
rect 127683 293147 127711 293175
rect 127497 293085 127525 293113
rect 127559 293085 127587 293113
rect 127621 293085 127649 293113
rect 127683 293085 127711 293113
rect 127497 293023 127525 293051
rect 127559 293023 127587 293051
rect 127621 293023 127649 293051
rect 127683 293023 127711 293051
rect 127497 292961 127525 292989
rect 127559 292961 127587 292989
rect 127621 292961 127649 292989
rect 127683 292961 127711 292989
rect 127497 284147 127525 284175
rect 127559 284147 127587 284175
rect 127621 284147 127649 284175
rect 127683 284147 127711 284175
rect 127497 284085 127525 284113
rect 127559 284085 127587 284113
rect 127621 284085 127649 284113
rect 127683 284085 127711 284113
rect 127497 284023 127525 284051
rect 127559 284023 127587 284051
rect 127621 284023 127649 284051
rect 127683 284023 127711 284051
rect 127497 283961 127525 283989
rect 127559 283961 127587 283989
rect 127621 283961 127649 283989
rect 127683 283961 127711 283989
rect 127497 275147 127525 275175
rect 127559 275147 127587 275175
rect 127621 275147 127649 275175
rect 127683 275147 127711 275175
rect 127497 275085 127525 275113
rect 127559 275085 127587 275113
rect 127621 275085 127649 275113
rect 127683 275085 127711 275113
rect 127497 275023 127525 275051
rect 127559 275023 127587 275051
rect 127621 275023 127649 275051
rect 127683 275023 127711 275051
rect 127497 274961 127525 274989
rect 127559 274961 127587 274989
rect 127621 274961 127649 274989
rect 127683 274961 127711 274989
rect 140997 298578 141025 298606
rect 141059 298578 141087 298606
rect 141121 298578 141149 298606
rect 141183 298578 141211 298606
rect 140997 298516 141025 298544
rect 141059 298516 141087 298544
rect 141121 298516 141149 298544
rect 141183 298516 141211 298544
rect 140997 298454 141025 298482
rect 141059 298454 141087 298482
rect 141121 298454 141149 298482
rect 141183 298454 141211 298482
rect 140997 298392 141025 298420
rect 141059 298392 141087 298420
rect 141121 298392 141149 298420
rect 141183 298392 141211 298420
rect 140997 290147 141025 290175
rect 141059 290147 141087 290175
rect 141121 290147 141149 290175
rect 141183 290147 141211 290175
rect 140997 290085 141025 290113
rect 141059 290085 141087 290113
rect 141121 290085 141149 290113
rect 141183 290085 141211 290113
rect 140997 290023 141025 290051
rect 141059 290023 141087 290051
rect 141121 290023 141149 290051
rect 141183 290023 141211 290051
rect 140997 289961 141025 289989
rect 141059 289961 141087 289989
rect 141121 289961 141149 289989
rect 141183 289961 141211 289989
rect 140997 281147 141025 281175
rect 141059 281147 141087 281175
rect 141121 281147 141149 281175
rect 141183 281147 141211 281175
rect 140997 281085 141025 281113
rect 141059 281085 141087 281113
rect 141121 281085 141149 281113
rect 141183 281085 141211 281113
rect 140997 281023 141025 281051
rect 141059 281023 141087 281051
rect 141121 281023 141149 281051
rect 141183 281023 141211 281051
rect 140997 280961 141025 280989
rect 141059 280961 141087 280989
rect 141121 280961 141149 280989
rect 141183 280961 141211 280989
rect 140997 272147 141025 272175
rect 141059 272147 141087 272175
rect 141121 272147 141149 272175
rect 141183 272147 141211 272175
rect 140997 272085 141025 272113
rect 141059 272085 141087 272113
rect 141121 272085 141149 272113
rect 141183 272085 141211 272113
rect 140997 272023 141025 272051
rect 141059 272023 141087 272051
rect 141121 272023 141149 272051
rect 141183 272023 141211 272051
rect 140997 271961 141025 271989
rect 141059 271961 141087 271989
rect 141121 271961 141149 271989
rect 141183 271961 141211 271989
rect 142857 299058 142885 299086
rect 142919 299058 142947 299086
rect 142981 299058 143009 299086
rect 143043 299058 143071 299086
rect 142857 298996 142885 299024
rect 142919 298996 142947 299024
rect 142981 298996 143009 299024
rect 143043 298996 143071 299024
rect 142857 298934 142885 298962
rect 142919 298934 142947 298962
rect 142981 298934 143009 298962
rect 143043 298934 143071 298962
rect 142857 298872 142885 298900
rect 142919 298872 142947 298900
rect 142981 298872 143009 298900
rect 143043 298872 143071 298900
rect 142857 293147 142885 293175
rect 142919 293147 142947 293175
rect 142981 293147 143009 293175
rect 143043 293147 143071 293175
rect 142857 293085 142885 293113
rect 142919 293085 142947 293113
rect 142981 293085 143009 293113
rect 143043 293085 143071 293113
rect 142857 293023 142885 293051
rect 142919 293023 142947 293051
rect 142981 293023 143009 293051
rect 143043 293023 143071 293051
rect 142857 292961 142885 292989
rect 142919 292961 142947 292989
rect 142981 292961 143009 292989
rect 143043 292961 143071 292989
rect 142857 284147 142885 284175
rect 142919 284147 142947 284175
rect 142981 284147 143009 284175
rect 143043 284147 143071 284175
rect 142857 284085 142885 284113
rect 142919 284085 142947 284113
rect 142981 284085 143009 284113
rect 143043 284085 143071 284113
rect 142857 284023 142885 284051
rect 142919 284023 142947 284051
rect 142981 284023 143009 284051
rect 143043 284023 143071 284051
rect 142857 283961 142885 283989
rect 142919 283961 142947 283989
rect 142981 283961 143009 283989
rect 143043 283961 143071 283989
rect 142857 275147 142885 275175
rect 142919 275147 142947 275175
rect 142981 275147 143009 275175
rect 143043 275147 143071 275175
rect 142857 275085 142885 275113
rect 142919 275085 142947 275113
rect 142981 275085 143009 275113
rect 143043 275085 143071 275113
rect 142857 275023 142885 275051
rect 142919 275023 142947 275051
rect 142981 275023 143009 275051
rect 143043 275023 143071 275051
rect 142857 274961 142885 274989
rect 142919 274961 142947 274989
rect 142981 274961 143009 274989
rect 143043 274961 143071 274989
rect 156357 298578 156385 298606
rect 156419 298578 156447 298606
rect 156481 298578 156509 298606
rect 156543 298578 156571 298606
rect 156357 298516 156385 298544
rect 156419 298516 156447 298544
rect 156481 298516 156509 298544
rect 156543 298516 156571 298544
rect 156357 298454 156385 298482
rect 156419 298454 156447 298482
rect 156481 298454 156509 298482
rect 156543 298454 156571 298482
rect 156357 298392 156385 298420
rect 156419 298392 156447 298420
rect 156481 298392 156509 298420
rect 156543 298392 156571 298420
rect 156357 290147 156385 290175
rect 156419 290147 156447 290175
rect 156481 290147 156509 290175
rect 156543 290147 156571 290175
rect 156357 290085 156385 290113
rect 156419 290085 156447 290113
rect 156481 290085 156509 290113
rect 156543 290085 156571 290113
rect 156357 290023 156385 290051
rect 156419 290023 156447 290051
rect 156481 290023 156509 290051
rect 156543 290023 156571 290051
rect 156357 289961 156385 289989
rect 156419 289961 156447 289989
rect 156481 289961 156509 289989
rect 156543 289961 156571 289989
rect 156357 281147 156385 281175
rect 156419 281147 156447 281175
rect 156481 281147 156509 281175
rect 156543 281147 156571 281175
rect 156357 281085 156385 281113
rect 156419 281085 156447 281113
rect 156481 281085 156509 281113
rect 156543 281085 156571 281113
rect 156357 281023 156385 281051
rect 156419 281023 156447 281051
rect 156481 281023 156509 281051
rect 156543 281023 156571 281051
rect 156357 280961 156385 280989
rect 156419 280961 156447 280989
rect 156481 280961 156509 280989
rect 156543 280961 156571 280989
rect 156357 272147 156385 272175
rect 156419 272147 156447 272175
rect 156481 272147 156509 272175
rect 156543 272147 156571 272175
rect 156357 272085 156385 272113
rect 156419 272085 156447 272113
rect 156481 272085 156509 272113
rect 156543 272085 156571 272113
rect 156357 272023 156385 272051
rect 156419 272023 156447 272051
rect 156481 272023 156509 272051
rect 156543 272023 156571 272051
rect 156357 271961 156385 271989
rect 156419 271961 156447 271989
rect 156481 271961 156509 271989
rect 156543 271961 156571 271989
rect 158217 299058 158245 299086
rect 158279 299058 158307 299086
rect 158341 299058 158369 299086
rect 158403 299058 158431 299086
rect 158217 298996 158245 299024
rect 158279 298996 158307 299024
rect 158341 298996 158369 299024
rect 158403 298996 158431 299024
rect 158217 298934 158245 298962
rect 158279 298934 158307 298962
rect 158341 298934 158369 298962
rect 158403 298934 158431 298962
rect 158217 298872 158245 298900
rect 158279 298872 158307 298900
rect 158341 298872 158369 298900
rect 158403 298872 158431 298900
rect 158217 293147 158245 293175
rect 158279 293147 158307 293175
rect 158341 293147 158369 293175
rect 158403 293147 158431 293175
rect 158217 293085 158245 293113
rect 158279 293085 158307 293113
rect 158341 293085 158369 293113
rect 158403 293085 158431 293113
rect 158217 293023 158245 293051
rect 158279 293023 158307 293051
rect 158341 293023 158369 293051
rect 158403 293023 158431 293051
rect 158217 292961 158245 292989
rect 158279 292961 158307 292989
rect 158341 292961 158369 292989
rect 158403 292961 158431 292989
rect 158217 284147 158245 284175
rect 158279 284147 158307 284175
rect 158341 284147 158369 284175
rect 158403 284147 158431 284175
rect 158217 284085 158245 284113
rect 158279 284085 158307 284113
rect 158341 284085 158369 284113
rect 158403 284085 158431 284113
rect 158217 284023 158245 284051
rect 158279 284023 158307 284051
rect 158341 284023 158369 284051
rect 158403 284023 158431 284051
rect 158217 283961 158245 283989
rect 158279 283961 158307 283989
rect 158341 283961 158369 283989
rect 158403 283961 158431 283989
rect 158217 275147 158245 275175
rect 158279 275147 158307 275175
rect 158341 275147 158369 275175
rect 158403 275147 158431 275175
rect 158217 275085 158245 275113
rect 158279 275085 158307 275113
rect 158341 275085 158369 275113
rect 158403 275085 158431 275113
rect 158217 275023 158245 275051
rect 158279 275023 158307 275051
rect 158341 275023 158369 275051
rect 158403 275023 158431 275051
rect 158217 274961 158245 274989
rect 158279 274961 158307 274989
rect 158341 274961 158369 274989
rect 158403 274961 158431 274989
rect 171717 298578 171745 298606
rect 171779 298578 171807 298606
rect 171841 298578 171869 298606
rect 171903 298578 171931 298606
rect 171717 298516 171745 298544
rect 171779 298516 171807 298544
rect 171841 298516 171869 298544
rect 171903 298516 171931 298544
rect 171717 298454 171745 298482
rect 171779 298454 171807 298482
rect 171841 298454 171869 298482
rect 171903 298454 171931 298482
rect 171717 298392 171745 298420
rect 171779 298392 171807 298420
rect 171841 298392 171869 298420
rect 171903 298392 171931 298420
rect 171717 290147 171745 290175
rect 171779 290147 171807 290175
rect 171841 290147 171869 290175
rect 171903 290147 171931 290175
rect 171717 290085 171745 290113
rect 171779 290085 171807 290113
rect 171841 290085 171869 290113
rect 171903 290085 171931 290113
rect 171717 290023 171745 290051
rect 171779 290023 171807 290051
rect 171841 290023 171869 290051
rect 171903 290023 171931 290051
rect 171717 289961 171745 289989
rect 171779 289961 171807 289989
rect 171841 289961 171869 289989
rect 171903 289961 171931 289989
rect 171717 281147 171745 281175
rect 171779 281147 171807 281175
rect 171841 281147 171869 281175
rect 171903 281147 171931 281175
rect 171717 281085 171745 281113
rect 171779 281085 171807 281113
rect 171841 281085 171869 281113
rect 171903 281085 171931 281113
rect 171717 281023 171745 281051
rect 171779 281023 171807 281051
rect 171841 281023 171869 281051
rect 171903 281023 171931 281051
rect 171717 280961 171745 280989
rect 171779 280961 171807 280989
rect 171841 280961 171869 280989
rect 171903 280961 171931 280989
rect 171717 272147 171745 272175
rect 171779 272147 171807 272175
rect 171841 272147 171869 272175
rect 171903 272147 171931 272175
rect 171717 272085 171745 272113
rect 171779 272085 171807 272113
rect 171841 272085 171869 272113
rect 171903 272085 171931 272113
rect 171717 272023 171745 272051
rect 171779 272023 171807 272051
rect 171841 272023 171869 272051
rect 171903 272023 171931 272051
rect 171717 271961 171745 271989
rect 171779 271961 171807 271989
rect 171841 271961 171869 271989
rect 171903 271961 171931 271989
rect 96777 266147 96805 266175
rect 96839 266147 96867 266175
rect 96901 266147 96929 266175
rect 96963 266147 96991 266175
rect 96777 266085 96805 266113
rect 96839 266085 96867 266113
rect 96901 266085 96929 266113
rect 96963 266085 96991 266113
rect 96777 266023 96805 266051
rect 96839 266023 96867 266051
rect 96901 266023 96929 266051
rect 96963 266023 96991 266051
rect 96777 265961 96805 265989
rect 96839 265961 96867 265989
rect 96901 265961 96929 265989
rect 96963 265961 96991 265989
rect 109939 266147 109967 266175
rect 110001 266147 110029 266175
rect 109939 266085 109967 266113
rect 110001 266085 110029 266113
rect 109939 266023 109967 266051
rect 110001 266023 110029 266051
rect 109939 265961 109967 265989
rect 110001 265961 110029 265989
rect 125299 266147 125327 266175
rect 125361 266147 125389 266175
rect 125299 266085 125327 266113
rect 125361 266085 125389 266113
rect 125299 266023 125327 266051
rect 125361 266023 125389 266051
rect 125299 265961 125327 265989
rect 125361 265961 125389 265989
rect 140659 266147 140687 266175
rect 140721 266147 140749 266175
rect 140659 266085 140687 266113
rect 140721 266085 140749 266113
rect 140659 266023 140687 266051
rect 140721 266023 140749 266051
rect 140659 265961 140687 265989
rect 140721 265961 140749 265989
rect 156019 266147 156047 266175
rect 156081 266147 156109 266175
rect 156019 266085 156047 266113
rect 156081 266085 156109 266113
rect 156019 266023 156047 266051
rect 156081 266023 156109 266051
rect 156019 265961 156047 265989
rect 156081 265961 156109 265989
rect 102259 263147 102287 263175
rect 102321 263147 102349 263175
rect 102259 263085 102287 263113
rect 102321 263085 102349 263113
rect 102259 263023 102287 263051
rect 102321 263023 102349 263051
rect 102259 262961 102287 262989
rect 102321 262961 102349 262989
rect 117619 263147 117647 263175
rect 117681 263147 117709 263175
rect 117619 263085 117647 263113
rect 117681 263085 117709 263113
rect 117619 263023 117647 263051
rect 117681 263023 117709 263051
rect 117619 262961 117647 262989
rect 117681 262961 117709 262989
rect 132979 263147 133007 263175
rect 133041 263147 133069 263175
rect 132979 263085 133007 263113
rect 133041 263085 133069 263113
rect 132979 263023 133007 263051
rect 133041 263023 133069 263051
rect 132979 262961 133007 262989
rect 133041 262961 133069 262989
rect 148339 263147 148367 263175
rect 148401 263147 148429 263175
rect 148339 263085 148367 263113
rect 148401 263085 148429 263113
rect 148339 263023 148367 263051
rect 148401 263023 148429 263051
rect 148339 262961 148367 262989
rect 148401 262961 148429 262989
rect 163699 263147 163727 263175
rect 163761 263147 163789 263175
rect 163699 263085 163727 263113
rect 163761 263085 163789 263113
rect 163699 263023 163727 263051
rect 163761 263023 163789 263051
rect 163699 262961 163727 262989
rect 163761 262961 163789 262989
rect 171717 263147 171745 263175
rect 171779 263147 171807 263175
rect 171841 263147 171869 263175
rect 171903 263147 171931 263175
rect 171717 263085 171745 263113
rect 171779 263085 171807 263113
rect 171841 263085 171869 263113
rect 171903 263085 171931 263113
rect 171717 263023 171745 263051
rect 171779 263023 171807 263051
rect 171841 263023 171869 263051
rect 171903 263023 171931 263051
rect 171717 262961 171745 262989
rect 171779 262961 171807 262989
rect 171841 262961 171869 262989
rect 171903 262961 171931 262989
rect 96777 257147 96805 257175
rect 96839 257147 96867 257175
rect 96901 257147 96929 257175
rect 96963 257147 96991 257175
rect 96777 257085 96805 257113
rect 96839 257085 96867 257113
rect 96901 257085 96929 257113
rect 96963 257085 96991 257113
rect 96777 257023 96805 257051
rect 96839 257023 96867 257051
rect 96901 257023 96929 257051
rect 96963 257023 96991 257051
rect 96777 256961 96805 256989
rect 96839 256961 96867 256989
rect 96901 256961 96929 256989
rect 96963 256961 96991 256989
rect 109939 257147 109967 257175
rect 110001 257147 110029 257175
rect 109939 257085 109967 257113
rect 110001 257085 110029 257113
rect 109939 257023 109967 257051
rect 110001 257023 110029 257051
rect 109939 256961 109967 256989
rect 110001 256961 110029 256989
rect 125299 257147 125327 257175
rect 125361 257147 125389 257175
rect 125299 257085 125327 257113
rect 125361 257085 125389 257113
rect 125299 257023 125327 257051
rect 125361 257023 125389 257051
rect 125299 256961 125327 256989
rect 125361 256961 125389 256989
rect 140659 257147 140687 257175
rect 140721 257147 140749 257175
rect 140659 257085 140687 257113
rect 140721 257085 140749 257113
rect 140659 257023 140687 257051
rect 140721 257023 140749 257051
rect 140659 256961 140687 256989
rect 140721 256961 140749 256989
rect 156019 257147 156047 257175
rect 156081 257147 156109 257175
rect 156019 257085 156047 257113
rect 156081 257085 156109 257113
rect 156019 257023 156047 257051
rect 156081 257023 156109 257051
rect 156019 256961 156047 256989
rect 156081 256961 156109 256989
rect 102259 254147 102287 254175
rect 102321 254147 102349 254175
rect 102259 254085 102287 254113
rect 102321 254085 102349 254113
rect 102259 254023 102287 254051
rect 102321 254023 102349 254051
rect 102259 253961 102287 253989
rect 102321 253961 102349 253989
rect 117619 254147 117647 254175
rect 117681 254147 117709 254175
rect 117619 254085 117647 254113
rect 117681 254085 117709 254113
rect 117619 254023 117647 254051
rect 117681 254023 117709 254051
rect 117619 253961 117647 253989
rect 117681 253961 117709 253989
rect 132979 254147 133007 254175
rect 133041 254147 133069 254175
rect 132979 254085 133007 254113
rect 133041 254085 133069 254113
rect 132979 254023 133007 254051
rect 133041 254023 133069 254051
rect 132979 253961 133007 253989
rect 133041 253961 133069 253989
rect 148339 254147 148367 254175
rect 148401 254147 148429 254175
rect 148339 254085 148367 254113
rect 148401 254085 148429 254113
rect 148339 254023 148367 254051
rect 148401 254023 148429 254051
rect 148339 253961 148367 253989
rect 148401 253961 148429 253989
rect 163699 254147 163727 254175
rect 163761 254147 163789 254175
rect 163699 254085 163727 254113
rect 163761 254085 163789 254113
rect 163699 254023 163727 254051
rect 163761 254023 163789 254051
rect 163699 253961 163727 253989
rect 163761 253961 163789 253989
rect 171717 254147 171745 254175
rect 171779 254147 171807 254175
rect 171841 254147 171869 254175
rect 171903 254147 171931 254175
rect 171717 254085 171745 254113
rect 171779 254085 171807 254113
rect 171841 254085 171869 254113
rect 171903 254085 171931 254113
rect 171717 254023 171745 254051
rect 171779 254023 171807 254051
rect 171841 254023 171869 254051
rect 171903 254023 171931 254051
rect 171717 253961 171745 253989
rect 171779 253961 171807 253989
rect 171841 253961 171869 253989
rect 171903 253961 171931 253989
rect 96777 248147 96805 248175
rect 96839 248147 96867 248175
rect 96901 248147 96929 248175
rect 96963 248147 96991 248175
rect 96777 248085 96805 248113
rect 96839 248085 96867 248113
rect 96901 248085 96929 248113
rect 96963 248085 96991 248113
rect 96777 248023 96805 248051
rect 96839 248023 96867 248051
rect 96901 248023 96929 248051
rect 96963 248023 96991 248051
rect 96777 247961 96805 247989
rect 96839 247961 96867 247989
rect 96901 247961 96929 247989
rect 96963 247961 96991 247989
rect 109939 248147 109967 248175
rect 110001 248147 110029 248175
rect 109939 248085 109967 248113
rect 110001 248085 110029 248113
rect 109939 248023 109967 248051
rect 110001 248023 110029 248051
rect 109939 247961 109967 247989
rect 110001 247961 110029 247989
rect 125299 248147 125327 248175
rect 125361 248147 125389 248175
rect 125299 248085 125327 248113
rect 125361 248085 125389 248113
rect 125299 248023 125327 248051
rect 125361 248023 125389 248051
rect 125299 247961 125327 247989
rect 125361 247961 125389 247989
rect 140659 248147 140687 248175
rect 140721 248147 140749 248175
rect 140659 248085 140687 248113
rect 140721 248085 140749 248113
rect 140659 248023 140687 248051
rect 140721 248023 140749 248051
rect 140659 247961 140687 247989
rect 140721 247961 140749 247989
rect 156019 248147 156047 248175
rect 156081 248147 156109 248175
rect 156019 248085 156047 248113
rect 156081 248085 156109 248113
rect 156019 248023 156047 248051
rect 156081 248023 156109 248051
rect 156019 247961 156047 247989
rect 156081 247961 156109 247989
rect 102259 245147 102287 245175
rect 102321 245147 102349 245175
rect 102259 245085 102287 245113
rect 102321 245085 102349 245113
rect 102259 245023 102287 245051
rect 102321 245023 102349 245051
rect 102259 244961 102287 244989
rect 102321 244961 102349 244989
rect 117619 245147 117647 245175
rect 117681 245147 117709 245175
rect 117619 245085 117647 245113
rect 117681 245085 117709 245113
rect 117619 245023 117647 245051
rect 117681 245023 117709 245051
rect 117619 244961 117647 244989
rect 117681 244961 117709 244989
rect 132979 245147 133007 245175
rect 133041 245147 133069 245175
rect 132979 245085 133007 245113
rect 133041 245085 133069 245113
rect 132979 245023 133007 245051
rect 133041 245023 133069 245051
rect 132979 244961 133007 244989
rect 133041 244961 133069 244989
rect 148339 245147 148367 245175
rect 148401 245147 148429 245175
rect 148339 245085 148367 245113
rect 148401 245085 148429 245113
rect 148339 245023 148367 245051
rect 148401 245023 148429 245051
rect 148339 244961 148367 244989
rect 148401 244961 148429 244989
rect 163699 245147 163727 245175
rect 163761 245147 163789 245175
rect 163699 245085 163727 245113
rect 163761 245085 163789 245113
rect 163699 245023 163727 245051
rect 163761 245023 163789 245051
rect 163699 244961 163727 244989
rect 163761 244961 163789 244989
rect 171717 245147 171745 245175
rect 171779 245147 171807 245175
rect 171841 245147 171869 245175
rect 171903 245147 171931 245175
rect 171717 245085 171745 245113
rect 171779 245085 171807 245113
rect 171841 245085 171869 245113
rect 171903 245085 171931 245113
rect 171717 245023 171745 245051
rect 171779 245023 171807 245051
rect 171841 245023 171869 245051
rect 171903 245023 171931 245051
rect 171717 244961 171745 244989
rect 171779 244961 171807 244989
rect 171841 244961 171869 244989
rect 171903 244961 171931 244989
rect 96777 239147 96805 239175
rect 96839 239147 96867 239175
rect 96901 239147 96929 239175
rect 96963 239147 96991 239175
rect 96777 239085 96805 239113
rect 96839 239085 96867 239113
rect 96901 239085 96929 239113
rect 96963 239085 96991 239113
rect 96777 239023 96805 239051
rect 96839 239023 96867 239051
rect 96901 239023 96929 239051
rect 96963 239023 96991 239051
rect 96777 238961 96805 238989
rect 96839 238961 96867 238989
rect 96901 238961 96929 238989
rect 96963 238961 96991 238989
rect 109939 239147 109967 239175
rect 110001 239147 110029 239175
rect 109939 239085 109967 239113
rect 110001 239085 110029 239113
rect 109939 239023 109967 239051
rect 110001 239023 110029 239051
rect 109939 238961 109967 238989
rect 110001 238961 110029 238989
rect 125299 239147 125327 239175
rect 125361 239147 125389 239175
rect 125299 239085 125327 239113
rect 125361 239085 125389 239113
rect 125299 239023 125327 239051
rect 125361 239023 125389 239051
rect 125299 238961 125327 238989
rect 125361 238961 125389 238989
rect 140659 239147 140687 239175
rect 140721 239147 140749 239175
rect 140659 239085 140687 239113
rect 140721 239085 140749 239113
rect 140659 239023 140687 239051
rect 140721 239023 140749 239051
rect 140659 238961 140687 238989
rect 140721 238961 140749 238989
rect 156019 239147 156047 239175
rect 156081 239147 156109 239175
rect 156019 239085 156047 239113
rect 156081 239085 156109 239113
rect 156019 239023 156047 239051
rect 156081 239023 156109 239051
rect 156019 238961 156047 238989
rect 156081 238961 156109 238989
rect 102259 236147 102287 236175
rect 102321 236147 102349 236175
rect 102259 236085 102287 236113
rect 102321 236085 102349 236113
rect 102259 236023 102287 236051
rect 102321 236023 102349 236051
rect 102259 235961 102287 235989
rect 102321 235961 102349 235989
rect 117619 236147 117647 236175
rect 117681 236147 117709 236175
rect 117619 236085 117647 236113
rect 117681 236085 117709 236113
rect 117619 236023 117647 236051
rect 117681 236023 117709 236051
rect 117619 235961 117647 235989
rect 117681 235961 117709 235989
rect 132979 236147 133007 236175
rect 133041 236147 133069 236175
rect 132979 236085 133007 236113
rect 133041 236085 133069 236113
rect 132979 236023 133007 236051
rect 133041 236023 133069 236051
rect 132979 235961 133007 235989
rect 133041 235961 133069 235989
rect 148339 236147 148367 236175
rect 148401 236147 148429 236175
rect 148339 236085 148367 236113
rect 148401 236085 148429 236113
rect 148339 236023 148367 236051
rect 148401 236023 148429 236051
rect 148339 235961 148367 235989
rect 148401 235961 148429 235989
rect 163699 236147 163727 236175
rect 163761 236147 163789 236175
rect 163699 236085 163727 236113
rect 163761 236085 163789 236113
rect 163699 236023 163727 236051
rect 163761 236023 163789 236051
rect 163699 235961 163727 235989
rect 163761 235961 163789 235989
rect 171717 236147 171745 236175
rect 171779 236147 171807 236175
rect 171841 236147 171869 236175
rect 171903 236147 171931 236175
rect 171717 236085 171745 236113
rect 171779 236085 171807 236113
rect 171841 236085 171869 236113
rect 171903 236085 171931 236113
rect 171717 236023 171745 236051
rect 171779 236023 171807 236051
rect 171841 236023 171869 236051
rect 171903 236023 171931 236051
rect 171717 235961 171745 235989
rect 171779 235961 171807 235989
rect 171841 235961 171869 235989
rect 171903 235961 171931 235989
rect 96777 230147 96805 230175
rect 96839 230147 96867 230175
rect 96901 230147 96929 230175
rect 96963 230147 96991 230175
rect 96777 230085 96805 230113
rect 96839 230085 96867 230113
rect 96901 230085 96929 230113
rect 96963 230085 96991 230113
rect 96777 230023 96805 230051
rect 96839 230023 96867 230051
rect 96901 230023 96929 230051
rect 96963 230023 96991 230051
rect 96777 229961 96805 229989
rect 96839 229961 96867 229989
rect 96901 229961 96929 229989
rect 96963 229961 96991 229989
rect 109939 230147 109967 230175
rect 110001 230147 110029 230175
rect 109939 230085 109967 230113
rect 110001 230085 110029 230113
rect 109939 230023 109967 230051
rect 110001 230023 110029 230051
rect 109939 229961 109967 229989
rect 110001 229961 110029 229989
rect 125299 230147 125327 230175
rect 125361 230147 125389 230175
rect 125299 230085 125327 230113
rect 125361 230085 125389 230113
rect 125299 230023 125327 230051
rect 125361 230023 125389 230051
rect 125299 229961 125327 229989
rect 125361 229961 125389 229989
rect 140659 230147 140687 230175
rect 140721 230147 140749 230175
rect 140659 230085 140687 230113
rect 140721 230085 140749 230113
rect 140659 230023 140687 230051
rect 140721 230023 140749 230051
rect 140659 229961 140687 229989
rect 140721 229961 140749 229989
rect 156019 230147 156047 230175
rect 156081 230147 156109 230175
rect 156019 230085 156047 230113
rect 156081 230085 156109 230113
rect 156019 230023 156047 230051
rect 156081 230023 156109 230051
rect 156019 229961 156047 229989
rect 156081 229961 156109 229989
rect 102259 227147 102287 227175
rect 102321 227147 102349 227175
rect 102259 227085 102287 227113
rect 102321 227085 102349 227113
rect 102259 227023 102287 227051
rect 102321 227023 102349 227051
rect 102259 226961 102287 226989
rect 102321 226961 102349 226989
rect 117619 227147 117647 227175
rect 117681 227147 117709 227175
rect 117619 227085 117647 227113
rect 117681 227085 117709 227113
rect 117619 227023 117647 227051
rect 117681 227023 117709 227051
rect 117619 226961 117647 226989
rect 117681 226961 117709 226989
rect 132979 227147 133007 227175
rect 133041 227147 133069 227175
rect 132979 227085 133007 227113
rect 133041 227085 133069 227113
rect 132979 227023 133007 227051
rect 133041 227023 133069 227051
rect 132979 226961 133007 226989
rect 133041 226961 133069 226989
rect 148339 227147 148367 227175
rect 148401 227147 148429 227175
rect 148339 227085 148367 227113
rect 148401 227085 148429 227113
rect 148339 227023 148367 227051
rect 148401 227023 148429 227051
rect 148339 226961 148367 226989
rect 148401 226961 148429 226989
rect 163699 227147 163727 227175
rect 163761 227147 163789 227175
rect 163699 227085 163727 227113
rect 163761 227085 163789 227113
rect 163699 227023 163727 227051
rect 163761 227023 163789 227051
rect 163699 226961 163727 226989
rect 163761 226961 163789 226989
rect 171717 227147 171745 227175
rect 171779 227147 171807 227175
rect 171841 227147 171869 227175
rect 171903 227147 171931 227175
rect 171717 227085 171745 227113
rect 171779 227085 171807 227113
rect 171841 227085 171869 227113
rect 171903 227085 171931 227113
rect 171717 227023 171745 227051
rect 171779 227023 171807 227051
rect 171841 227023 171869 227051
rect 171903 227023 171931 227051
rect 171717 226961 171745 226989
rect 171779 226961 171807 226989
rect 171841 226961 171869 226989
rect 171903 226961 171931 226989
rect 96777 221147 96805 221175
rect 96839 221147 96867 221175
rect 96901 221147 96929 221175
rect 96963 221147 96991 221175
rect 96777 221085 96805 221113
rect 96839 221085 96867 221113
rect 96901 221085 96929 221113
rect 96963 221085 96991 221113
rect 96777 221023 96805 221051
rect 96839 221023 96867 221051
rect 96901 221023 96929 221051
rect 96963 221023 96991 221051
rect 96777 220961 96805 220989
rect 96839 220961 96867 220989
rect 96901 220961 96929 220989
rect 96963 220961 96991 220989
rect 109939 221147 109967 221175
rect 110001 221147 110029 221175
rect 109939 221085 109967 221113
rect 110001 221085 110029 221113
rect 109939 221023 109967 221051
rect 110001 221023 110029 221051
rect 109939 220961 109967 220989
rect 110001 220961 110029 220989
rect 125299 221147 125327 221175
rect 125361 221147 125389 221175
rect 125299 221085 125327 221113
rect 125361 221085 125389 221113
rect 125299 221023 125327 221051
rect 125361 221023 125389 221051
rect 125299 220961 125327 220989
rect 125361 220961 125389 220989
rect 140659 221147 140687 221175
rect 140721 221147 140749 221175
rect 140659 221085 140687 221113
rect 140721 221085 140749 221113
rect 140659 221023 140687 221051
rect 140721 221023 140749 221051
rect 140659 220961 140687 220989
rect 140721 220961 140749 220989
rect 156019 221147 156047 221175
rect 156081 221147 156109 221175
rect 156019 221085 156047 221113
rect 156081 221085 156109 221113
rect 156019 221023 156047 221051
rect 156081 221023 156109 221051
rect 156019 220961 156047 220989
rect 156081 220961 156109 220989
rect 102259 218147 102287 218175
rect 102321 218147 102349 218175
rect 102259 218085 102287 218113
rect 102321 218085 102349 218113
rect 102259 218023 102287 218051
rect 102321 218023 102349 218051
rect 102259 217961 102287 217989
rect 102321 217961 102349 217989
rect 117619 218147 117647 218175
rect 117681 218147 117709 218175
rect 117619 218085 117647 218113
rect 117681 218085 117709 218113
rect 117619 218023 117647 218051
rect 117681 218023 117709 218051
rect 117619 217961 117647 217989
rect 117681 217961 117709 217989
rect 132979 218147 133007 218175
rect 133041 218147 133069 218175
rect 132979 218085 133007 218113
rect 133041 218085 133069 218113
rect 132979 218023 133007 218051
rect 133041 218023 133069 218051
rect 132979 217961 133007 217989
rect 133041 217961 133069 217989
rect 148339 218147 148367 218175
rect 148401 218147 148429 218175
rect 148339 218085 148367 218113
rect 148401 218085 148429 218113
rect 148339 218023 148367 218051
rect 148401 218023 148429 218051
rect 148339 217961 148367 217989
rect 148401 217961 148429 217989
rect 163699 218147 163727 218175
rect 163761 218147 163789 218175
rect 163699 218085 163727 218113
rect 163761 218085 163789 218113
rect 163699 218023 163727 218051
rect 163761 218023 163789 218051
rect 163699 217961 163727 217989
rect 163761 217961 163789 217989
rect 171717 218147 171745 218175
rect 171779 218147 171807 218175
rect 171841 218147 171869 218175
rect 171903 218147 171931 218175
rect 171717 218085 171745 218113
rect 171779 218085 171807 218113
rect 171841 218085 171869 218113
rect 171903 218085 171931 218113
rect 171717 218023 171745 218051
rect 171779 218023 171807 218051
rect 171841 218023 171869 218051
rect 171903 218023 171931 218051
rect 171717 217961 171745 217989
rect 171779 217961 171807 217989
rect 171841 217961 171869 217989
rect 171903 217961 171931 217989
rect 96777 212147 96805 212175
rect 96839 212147 96867 212175
rect 96901 212147 96929 212175
rect 96963 212147 96991 212175
rect 96777 212085 96805 212113
rect 96839 212085 96867 212113
rect 96901 212085 96929 212113
rect 96963 212085 96991 212113
rect 96777 212023 96805 212051
rect 96839 212023 96867 212051
rect 96901 212023 96929 212051
rect 96963 212023 96991 212051
rect 96777 211961 96805 211989
rect 96839 211961 96867 211989
rect 96901 211961 96929 211989
rect 96963 211961 96991 211989
rect 109939 212147 109967 212175
rect 110001 212147 110029 212175
rect 109939 212085 109967 212113
rect 110001 212085 110029 212113
rect 109939 212023 109967 212051
rect 110001 212023 110029 212051
rect 109939 211961 109967 211989
rect 110001 211961 110029 211989
rect 125299 212147 125327 212175
rect 125361 212147 125389 212175
rect 125299 212085 125327 212113
rect 125361 212085 125389 212113
rect 125299 212023 125327 212051
rect 125361 212023 125389 212051
rect 125299 211961 125327 211989
rect 125361 211961 125389 211989
rect 140659 212147 140687 212175
rect 140721 212147 140749 212175
rect 140659 212085 140687 212113
rect 140721 212085 140749 212113
rect 140659 212023 140687 212051
rect 140721 212023 140749 212051
rect 140659 211961 140687 211989
rect 140721 211961 140749 211989
rect 156019 212147 156047 212175
rect 156081 212147 156109 212175
rect 156019 212085 156047 212113
rect 156081 212085 156109 212113
rect 156019 212023 156047 212051
rect 156081 212023 156109 212051
rect 156019 211961 156047 211989
rect 156081 211961 156109 211989
rect 102259 209147 102287 209175
rect 102321 209147 102349 209175
rect 102259 209085 102287 209113
rect 102321 209085 102349 209113
rect 102259 209023 102287 209051
rect 102321 209023 102349 209051
rect 102259 208961 102287 208989
rect 102321 208961 102349 208989
rect 117619 209147 117647 209175
rect 117681 209147 117709 209175
rect 117619 209085 117647 209113
rect 117681 209085 117709 209113
rect 117619 209023 117647 209051
rect 117681 209023 117709 209051
rect 117619 208961 117647 208989
rect 117681 208961 117709 208989
rect 132979 209147 133007 209175
rect 133041 209147 133069 209175
rect 132979 209085 133007 209113
rect 133041 209085 133069 209113
rect 132979 209023 133007 209051
rect 133041 209023 133069 209051
rect 132979 208961 133007 208989
rect 133041 208961 133069 208989
rect 148339 209147 148367 209175
rect 148401 209147 148429 209175
rect 148339 209085 148367 209113
rect 148401 209085 148429 209113
rect 148339 209023 148367 209051
rect 148401 209023 148429 209051
rect 148339 208961 148367 208989
rect 148401 208961 148429 208989
rect 163699 209147 163727 209175
rect 163761 209147 163789 209175
rect 163699 209085 163727 209113
rect 163761 209085 163789 209113
rect 163699 209023 163727 209051
rect 163761 209023 163789 209051
rect 163699 208961 163727 208989
rect 163761 208961 163789 208989
rect 171717 209147 171745 209175
rect 171779 209147 171807 209175
rect 171841 209147 171869 209175
rect 171903 209147 171931 209175
rect 171717 209085 171745 209113
rect 171779 209085 171807 209113
rect 171841 209085 171869 209113
rect 171903 209085 171931 209113
rect 171717 209023 171745 209051
rect 171779 209023 171807 209051
rect 171841 209023 171869 209051
rect 171903 209023 171931 209051
rect 171717 208961 171745 208989
rect 171779 208961 171807 208989
rect 171841 208961 171869 208989
rect 171903 208961 171931 208989
rect 96777 203147 96805 203175
rect 96839 203147 96867 203175
rect 96901 203147 96929 203175
rect 96963 203147 96991 203175
rect 96777 203085 96805 203113
rect 96839 203085 96867 203113
rect 96901 203085 96929 203113
rect 96963 203085 96991 203113
rect 96777 203023 96805 203051
rect 96839 203023 96867 203051
rect 96901 203023 96929 203051
rect 96963 203023 96991 203051
rect 96777 202961 96805 202989
rect 96839 202961 96867 202989
rect 96901 202961 96929 202989
rect 96963 202961 96991 202989
rect 109939 203147 109967 203175
rect 110001 203147 110029 203175
rect 109939 203085 109967 203113
rect 110001 203085 110029 203113
rect 109939 203023 109967 203051
rect 110001 203023 110029 203051
rect 109939 202961 109967 202989
rect 110001 202961 110029 202989
rect 125299 203147 125327 203175
rect 125361 203147 125389 203175
rect 125299 203085 125327 203113
rect 125361 203085 125389 203113
rect 125299 203023 125327 203051
rect 125361 203023 125389 203051
rect 125299 202961 125327 202989
rect 125361 202961 125389 202989
rect 140659 203147 140687 203175
rect 140721 203147 140749 203175
rect 140659 203085 140687 203113
rect 140721 203085 140749 203113
rect 140659 203023 140687 203051
rect 140721 203023 140749 203051
rect 140659 202961 140687 202989
rect 140721 202961 140749 202989
rect 156019 203147 156047 203175
rect 156081 203147 156109 203175
rect 156019 203085 156047 203113
rect 156081 203085 156109 203113
rect 156019 203023 156047 203051
rect 156081 203023 156109 203051
rect 156019 202961 156047 202989
rect 156081 202961 156109 202989
rect 102259 200147 102287 200175
rect 102321 200147 102349 200175
rect 102259 200085 102287 200113
rect 102321 200085 102349 200113
rect 102259 200023 102287 200051
rect 102321 200023 102349 200051
rect 102259 199961 102287 199989
rect 102321 199961 102349 199989
rect 117619 200147 117647 200175
rect 117681 200147 117709 200175
rect 117619 200085 117647 200113
rect 117681 200085 117709 200113
rect 117619 200023 117647 200051
rect 117681 200023 117709 200051
rect 117619 199961 117647 199989
rect 117681 199961 117709 199989
rect 132979 200147 133007 200175
rect 133041 200147 133069 200175
rect 132979 200085 133007 200113
rect 133041 200085 133069 200113
rect 132979 200023 133007 200051
rect 133041 200023 133069 200051
rect 132979 199961 133007 199989
rect 133041 199961 133069 199989
rect 148339 200147 148367 200175
rect 148401 200147 148429 200175
rect 148339 200085 148367 200113
rect 148401 200085 148429 200113
rect 148339 200023 148367 200051
rect 148401 200023 148429 200051
rect 148339 199961 148367 199989
rect 148401 199961 148429 199989
rect 163699 200147 163727 200175
rect 163761 200147 163789 200175
rect 163699 200085 163727 200113
rect 163761 200085 163789 200113
rect 163699 200023 163727 200051
rect 163761 200023 163789 200051
rect 163699 199961 163727 199989
rect 163761 199961 163789 199989
rect 171717 200147 171745 200175
rect 171779 200147 171807 200175
rect 171841 200147 171869 200175
rect 171903 200147 171931 200175
rect 171717 200085 171745 200113
rect 171779 200085 171807 200113
rect 171841 200085 171869 200113
rect 171903 200085 171931 200113
rect 171717 200023 171745 200051
rect 171779 200023 171807 200051
rect 171841 200023 171869 200051
rect 171903 200023 171931 200051
rect 171717 199961 171745 199989
rect 171779 199961 171807 199989
rect 171841 199961 171869 199989
rect 171903 199961 171931 199989
rect 96777 194147 96805 194175
rect 96839 194147 96867 194175
rect 96901 194147 96929 194175
rect 96963 194147 96991 194175
rect 96777 194085 96805 194113
rect 96839 194085 96867 194113
rect 96901 194085 96929 194113
rect 96963 194085 96991 194113
rect 96777 194023 96805 194051
rect 96839 194023 96867 194051
rect 96901 194023 96929 194051
rect 96963 194023 96991 194051
rect 96777 193961 96805 193989
rect 96839 193961 96867 193989
rect 96901 193961 96929 193989
rect 96963 193961 96991 193989
rect 109939 194147 109967 194175
rect 110001 194147 110029 194175
rect 109939 194085 109967 194113
rect 110001 194085 110029 194113
rect 109939 194023 109967 194051
rect 110001 194023 110029 194051
rect 109939 193961 109967 193989
rect 110001 193961 110029 193989
rect 125299 194147 125327 194175
rect 125361 194147 125389 194175
rect 125299 194085 125327 194113
rect 125361 194085 125389 194113
rect 125299 194023 125327 194051
rect 125361 194023 125389 194051
rect 125299 193961 125327 193989
rect 125361 193961 125389 193989
rect 140659 194147 140687 194175
rect 140721 194147 140749 194175
rect 140659 194085 140687 194113
rect 140721 194085 140749 194113
rect 140659 194023 140687 194051
rect 140721 194023 140749 194051
rect 140659 193961 140687 193989
rect 140721 193961 140749 193989
rect 156019 194147 156047 194175
rect 156081 194147 156109 194175
rect 156019 194085 156047 194113
rect 156081 194085 156109 194113
rect 156019 194023 156047 194051
rect 156081 194023 156109 194051
rect 156019 193961 156047 193989
rect 156081 193961 156109 193989
rect 102259 191147 102287 191175
rect 102321 191147 102349 191175
rect 102259 191085 102287 191113
rect 102321 191085 102349 191113
rect 102259 191023 102287 191051
rect 102321 191023 102349 191051
rect 102259 190961 102287 190989
rect 102321 190961 102349 190989
rect 117619 191147 117647 191175
rect 117681 191147 117709 191175
rect 117619 191085 117647 191113
rect 117681 191085 117709 191113
rect 117619 191023 117647 191051
rect 117681 191023 117709 191051
rect 117619 190961 117647 190989
rect 117681 190961 117709 190989
rect 132979 191147 133007 191175
rect 133041 191147 133069 191175
rect 132979 191085 133007 191113
rect 133041 191085 133069 191113
rect 132979 191023 133007 191051
rect 133041 191023 133069 191051
rect 132979 190961 133007 190989
rect 133041 190961 133069 190989
rect 148339 191147 148367 191175
rect 148401 191147 148429 191175
rect 148339 191085 148367 191113
rect 148401 191085 148429 191113
rect 148339 191023 148367 191051
rect 148401 191023 148429 191051
rect 148339 190961 148367 190989
rect 148401 190961 148429 190989
rect 163699 191147 163727 191175
rect 163761 191147 163789 191175
rect 163699 191085 163727 191113
rect 163761 191085 163789 191113
rect 163699 191023 163727 191051
rect 163761 191023 163789 191051
rect 163699 190961 163727 190989
rect 163761 190961 163789 190989
rect 171717 191147 171745 191175
rect 171779 191147 171807 191175
rect 171841 191147 171869 191175
rect 171903 191147 171931 191175
rect 171717 191085 171745 191113
rect 171779 191085 171807 191113
rect 171841 191085 171869 191113
rect 171903 191085 171931 191113
rect 171717 191023 171745 191051
rect 171779 191023 171807 191051
rect 171841 191023 171869 191051
rect 171903 191023 171931 191051
rect 171717 190961 171745 190989
rect 171779 190961 171807 190989
rect 171841 190961 171869 190989
rect 171903 190961 171931 190989
rect 96777 185147 96805 185175
rect 96839 185147 96867 185175
rect 96901 185147 96929 185175
rect 96963 185147 96991 185175
rect 96777 185085 96805 185113
rect 96839 185085 96867 185113
rect 96901 185085 96929 185113
rect 96963 185085 96991 185113
rect 96777 185023 96805 185051
rect 96839 185023 96867 185051
rect 96901 185023 96929 185051
rect 96963 185023 96991 185051
rect 96777 184961 96805 184989
rect 96839 184961 96867 184989
rect 96901 184961 96929 184989
rect 96963 184961 96991 184989
rect 109939 185147 109967 185175
rect 110001 185147 110029 185175
rect 109939 185085 109967 185113
rect 110001 185085 110029 185113
rect 109939 185023 109967 185051
rect 110001 185023 110029 185051
rect 109939 184961 109967 184989
rect 110001 184961 110029 184989
rect 125299 185147 125327 185175
rect 125361 185147 125389 185175
rect 125299 185085 125327 185113
rect 125361 185085 125389 185113
rect 125299 185023 125327 185051
rect 125361 185023 125389 185051
rect 125299 184961 125327 184989
rect 125361 184961 125389 184989
rect 140659 185147 140687 185175
rect 140721 185147 140749 185175
rect 140659 185085 140687 185113
rect 140721 185085 140749 185113
rect 140659 185023 140687 185051
rect 140721 185023 140749 185051
rect 140659 184961 140687 184989
rect 140721 184961 140749 184989
rect 156019 185147 156047 185175
rect 156081 185147 156109 185175
rect 156019 185085 156047 185113
rect 156081 185085 156109 185113
rect 156019 185023 156047 185051
rect 156081 185023 156109 185051
rect 156019 184961 156047 184989
rect 156081 184961 156109 184989
rect 102259 182147 102287 182175
rect 102321 182147 102349 182175
rect 102259 182085 102287 182113
rect 102321 182085 102349 182113
rect 102259 182023 102287 182051
rect 102321 182023 102349 182051
rect 102259 181961 102287 181989
rect 102321 181961 102349 181989
rect 117619 182147 117647 182175
rect 117681 182147 117709 182175
rect 117619 182085 117647 182113
rect 117681 182085 117709 182113
rect 117619 182023 117647 182051
rect 117681 182023 117709 182051
rect 117619 181961 117647 181989
rect 117681 181961 117709 181989
rect 132979 182147 133007 182175
rect 133041 182147 133069 182175
rect 132979 182085 133007 182113
rect 133041 182085 133069 182113
rect 132979 182023 133007 182051
rect 133041 182023 133069 182051
rect 132979 181961 133007 181989
rect 133041 181961 133069 181989
rect 148339 182147 148367 182175
rect 148401 182147 148429 182175
rect 148339 182085 148367 182113
rect 148401 182085 148429 182113
rect 148339 182023 148367 182051
rect 148401 182023 148429 182051
rect 148339 181961 148367 181989
rect 148401 181961 148429 181989
rect 163699 182147 163727 182175
rect 163761 182147 163789 182175
rect 163699 182085 163727 182113
rect 163761 182085 163789 182113
rect 163699 182023 163727 182051
rect 163761 182023 163789 182051
rect 163699 181961 163727 181989
rect 163761 181961 163789 181989
rect 171717 182147 171745 182175
rect 171779 182147 171807 182175
rect 171841 182147 171869 182175
rect 171903 182147 171931 182175
rect 171717 182085 171745 182113
rect 171779 182085 171807 182113
rect 171841 182085 171869 182113
rect 171903 182085 171931 182113
rect 171717 182023 171745 182051
rect 171779 182023 171807 182051
rect 171841 182023 171869 182051
rect 171903 182023 171931 182051
rect 171717 181961 171745 181989
rect 171779 181961 171807 181989
rect 171841 181961 171869 181989
rect 171903 181961 171931 181989
rect 96777 176147 96805 176175
rect 96839 176147 96867 176175
rect 96901 176147 96929 176175
rect 96963 176147 96991 176175
rect 96777 176085 96805 176113
rect 96839 176085 96867 176113
rect 96901 176085 96929 176113
rect 96963 176085 96991 176113
rect 96777 176023 96805 176051
rect 96839 176023 96867 176051
rect 96901 176023 96929 176051
rect 96963 176023 96991 176051
rect 96777 175961 96805 175989
rect 96839 175961 96867 175989
rect 96901 175961 96929 175989
rect 96963 175961 96991 175989
rect 109939 176147 109967 176175
rect 110001 176147 110029 176175
rect 109939 176085 109967 176113
rect 110001 176085 110029 176113
rect 109939 176023 109967 176051
rect 110001 176023 110029 176051
rect 109939 175961 109967 175989
rect 110001 175961 110029 175989
rect 125299 176147 125327 176175
rect 125361 176147 125389 176175
rect 125299 176085 125327 176113
rect 125361 176085 125389 176113
rect 125299 176023 125327 176051
rect 125361 176023 125389 176051
rect 125299 175961 125327 175989
rect 125361 175961 125389 175989
rect 140659 176147 140687 176175
rect 140721 176147 140749 176175
rect 140659 176085 140687 176113
rect 140721 176085 140749 176113
rect 140659 176023 140687 176051
rect 140721 176023 140749 176051
rect 140659 175961 140687 175989
rect 140721 175961 140749 175989
rect 156019 176147 156047 176175
rect 156081 176147 156109 176175
rect 156019 176085 156047 176113
rect 156081 176085 156109 176113
rect 156019 176023 156047 176051
rect 156081 176023 156109 176051
rect 156019 175961 156047 175989
rect 156081 175961 156109 175989
rect 102259 173147 102287 173175
rect 102321 173147 102349 173175
rect 102259 173085 102287 173113
rect 102321 173085 102349 173113
rect 102259 173023 102287 173051
rect 102321 173023 102349 173051
rect 102259 172961 102287 172989
rect 102321 172961 102349 172989
rect 117619 173147 117647 173175
rect 117681 173147 117709 173175
rect 117619 173085 117647 173113
rect 117681 173085 117709 173113
rect 117619 173023 117647 173051
rect 117681 173023 117709 173051
rect 117619 172961 117647 172989
rect 117681 172961 117709 172989
rect 132979 173147 133007 173175
rect 133041 173147 133069 173175
rect 132979 173085 133007 173113
rect 133041 173085 133069 173113
rect 132979 173023 133007 173051
rect 133041 173023 133069 173051
rect 132979 172961 133007 172989
rect 133041 172961 133069 172989
rect 148339 173147 148367 173175
rect 148401 173147 148429 173175
rect 148339 173085 148367 173113
rect 148401 173085 148429 173113
rect 148339 173023 148367 173051
rect 148401 173023 148429 173051
rect 148339 172961 148367 172989
rect 148401 172961 148429 172989
rect 163699 173147 163727 173175
rect 163761 173147 163789 173175
rect 163699 173085 163727 173113
rect 163761 173085 163789 173113
rect 163699 173023 163727 173051
rect 163761 173023 163789 173051
rect 163699 172961 163727 172989
rect 163761 172961 163789 172989
rect 171717 173147 171745 173175
rect 171779 173147 171807 173175
rect 171841 173147 171869 173175
rect 171903 173147 171931 173175
rect 171717 173085 171745 173113
rect 171779 173085 171807 173113
rect 171841 173085 171869 173113
rect 171903 173085 171931 173113
rect 171717 173023 171745 173051
rect 171779 173023 171807 173051
rect 171841 173023 171869 173051
rect 171903 173023 171931 173051
rect 171717 172961 171745 172989
rect 171779 172961 171807 172989
rect 171841 172961 171869 172989
rect 171903 172961 171931 172989
rect 96777 167147 96805 167175
rect 96839 167147 96867 167175
rect 96901 167147 96929 167175
rect 96963 167147 96991 167175
rect 96777 167085 96805 167113
rect 96839 167085 96867 167113
rect 96901 167085 96929 167113
rect 96963 167085 96991 167113
rect 96777 167023 96805 167051
rect 96839 167023 96867 167051
rect 96901 167023 96929 167051
rect 96963 167023 96991 167051
rect 96777 166961 96805 166989
rect 96839 166961 96867 166989
rect 96901 166961 96929 166989
rect 96963 166961 96991 166989
rect 171717 164147 171745 164175
rect 171779 164147 171807 164175
rect 171841 164147 171869 164175
rect 171903 164147 171931 164175
rect 171717 164085 171745 164113
rect 171779 164085 171807 164113
rect 171841 164085 171869 164113
rect 171903 164085 171931 164113
rect 171717 164023 171745 164051
rect 171779 164023 171807 164051
rect 171841 164023 171869 164051
rect 171903 164023 171931 164051
rect 171717 163961 171745 163989
rect 171779 163961 171807 163989
rect 171841 163961 171869 163989
rect 171903 163961 171931 163989
rect 173577 299058 173605 299086
rect 173639 299058 173667 299086
rect 173701 299058 173729 299086
rect 173763 299058 173791 299086
rect 173577 298996 173605 299024
rect 173639 298996 173667 299024
rect 173701 298996 173729 299024
rect 173763 298996 173791 299024
rect 173577 298934 173605 298962
rect 173639 298934 173667 298962
rect 173701 298934 173729 298962
rect 173763 298934 173791 298962
rect 173577 298872 173605 298900
rect 173639 298872 173667 298900
rect 173701 298872 173729 298900
rect 173763 298872 173791 298900
rect 173577 293147 173605 293175
rect 173639 293147 173667 293175
rect 173701 293147 173729 293175
rect 173763 293147 173791 293175
rect 173577 293085 173605 293113
rect 173639 293085 173667 293113
rect 173701 293085 173729 293113
rect 173763 293085 173791 293113
rect 173577 293023 173605 293051
rect 173639 293023 173667 293051
rect 173701 293023 173729 293051
rect 173763 293023 173791 293051
rect 173577 292961 173605 292989
rect 173639 292961 173667 292989
rect 173701 292961 173729 292989
rect 173763 292961 173791 292989
rect 173577 284147 173605 284175
rect 173639 284147 173667 284175
rect 173701 284147 173729 284175
rect 173763 284147 173791 284175
rect 173577 284085 173605 284113
rect 173639 284085 173667 284113
rect 173701 284085 173729 284113
rect 173763 284085 173791 284113
rect 173577 284023 173605 284051
rect 173639 284023 173667 284051
rect 173701 284023 173729 284051
rect 173763 284023 173791 284051
rect 173577 283961 173605 283989
rect 173639 283961 173667 283989
rect 173701 283961 173729 283989
rect 173763 283961 173791 283989
rect 173577 275147 173605 275175
rect 173639 275147 173667 275175
rect 173701 275147 173729 275175
rect 173763 275147 173791 275175
rect 173577 275085 173605 275113
rect 173639 275085 173667 275113
rect 173701 275085 173729 275113
rect 173763 275085 173791 275113
rect 173577 275023 173605 275051
rect 173639 275023 173667 275051
rect 173701 275023 173729 275051
rect 173763 275023 173791 275051
rect 173577 274961 173605 274989
rect 173639 274961 173667 274989
rect 173701 274961 173729 274989
rect 173763 274961 173791 274989
rect 173577 266147 173605 266175
rect 173639 266147 173667 266175
rect 173701 266147 173729 266175
rect 173763 266147 173791 266175
rect 173577 266085 173605 266113
rect 173639 266085 173667 266113
rect 173701 266085 173729 266113
rect 173763 266085 173791 266113
rect 173577 266023 173605 266051
rect 173639 266023 173667 266051
rect 173701 266023 173729 266051
rect 173763 266023 173791 266051
rect 173577 265961 173605 265989
rect 173639 265961 173667 265989
rect 173701 265961 173729 265989
rect 173763 265961 173791 265989
rect 173577 257147 173605 257175
rect 173639 257147 173667 257175
rect 173701 257147 173729 257175
rect 173763 257147 173791 257175
rect 173577 257085 173605 257113
rect 173639 257085 173667 257113
rect 173701 257085 173729 257113
rect 173763 257085 173791 257113
rect 173577 257023 173605 257051
rect 173639 257023 173667 257051
rect 173701 257023 173729 257051
rect 173763 257023 173791 257051
rect 173577 256961 173605 256989
rect 173639 256961 173667 256989
rect 173701 256961 173729 256989
rect 173763 256961 173791 256989
rect 173577 248147 173605 248175
rect 173639 248147 173667 248175
rect 173701 248147 173729 248175
rect 173763 248147 173791 248175
rect 173577 248085 173605 248113
rect 173639 248085 173667 248113
rect 173701 248085 173729 248113
rect 173763 248085 173791 248113
rect 173577 248023 173605 248051
rect 173639 248023 173667 248051
rect 173701 248023 173729 248051
rect 173763 248023 173791 248051
rect 173577 247961 173605 247989
rect 173639 247961 173667 247989
rect 173701 247961 173729 247989
rect 173763 247961 173791 247989
rect 173577 239147 173605 239175
rect 173639 239147 173667 239175
rect 173701 239147 173729 239175
rect 173763 239147 173791 239175
rect 173577 239085 173605 239113
rect 173639 239085 173667 239113
rect 173701 239085 173729 239113
rect 173763 239085 173791 239113
rect 173577 239023 173605 239051
rect 173639 239023 173667 239051
rect 173701 239023 173729 239051
rect 173763 239023 173791 239051
rect 173577 238961 173605 238989
rect 173639 238961 173667 238989
rect 173701 238961 173729 238989
rect 173763 238961 173791 238989
rect 173577 230147 173605 230175
rect 173639 230147 173667 230175
rect 173701 230147 173729 230175
rect 173763 230147 173791 230175
rect 173577 230085 173605 230113
rect 173639 230085 173667 230113
rect 173701 230085 173729 230113
rect 173763 230085 173791 230113
rect 173577 230023 173605 230051
rect 173639 230023 173667 230051
rect 173701 230023 173729 230051
rect 173763 230023 173791 230051
rect 173577 229961 173605 229989
rect 173639 229961 173667 229989
rect 173701 229961 173729 229989
rect 173763 229961 173791 229989
rect 173577 221147 173605 221175
rect 173639 221147 173667 221175
rect 173701 221147 173729 221175
rect 173763 221147 173791 221175
rect 173577 221085 173605 221113
rect 173639 221085 173667 221113
rect 173701 221085 173729 221113
rect 173763 221085 173791 221113
rect 173577 221023 173605 221051
rect 173639 221023 173667 221051
rect 173701 221023 173729 221051
rect 173763 221023 173791 221051
rect 173577 220961 173605 220989
rect 173639 220961 173667 220989
rect 173701 220961 173729 220989
rect 173763 220961 173791 220989
rect 173577 212147 173605 212175
rect 173639 212147 173667 212175
rect 173701 212147 173729 212175
rect 173763 212147 173791 212175
rect 173577 212085 173605 212113
rect 173639 212085 173667 212113
rect 173701 212085 173729 212113
rect 173763 212085 173791 212113
rect 173577 212023 173605 212051
rect 173639 212023 173667 212051
rect 173701 212023 173729 212051
rect 173763 212023 173791 212051
rect 173577 211961 173605 211989
rect 173639 211961 173667 211989
rect 173701 211961 173729 211989
rect 173763 211961 173791 211989
rect 173577 203147 173605 203175
rect 173639 203147 173667 203175
rect 173701 203147 173729 203175
rect 173763 203147 173791 203175
rect 173577 203085 173605 203113
rect 173639 203085 173667 203113
rect 173701 203085 173729 203113
rect 173763 203085 173791 203113
rect 173577 203023 173605 203051
rect 173639 203023 173667 203051
rect 173701 203023 173729 203051
rect 173763 203023 173791 203051
rect 173577 202961 173605 202989
rect 173639 202961 173667 202989
rect 173701 202961 173729 202989
rect 173763 202961 173791 202989
rect 173577 194147 173605 194175
rect 173639 194147 173667 194175
rect 173701 194147 173729 194175
rect 173763 194147 173791 194175
rect 173577 194085 173605 194113
rect 173639 194085 173667 194113
rect 173701 194085 173729 194113
rect 173763 194085 173791 194113
rect 173577 194023 173605 194051
rect 173639 194023 173667 194051
rect 173701 194023 173729 194051
rect 173763 194023 173791 194051
rect 173577 193961 173605 193989
rect 173639 193961 173667 193989
rect 173701 193961 173729 193989
rect 173763 193961 173791 193989
rect 187077 298578 187105 298606
rect 187139 298578 187167 298606
rect 187201 298578 187229 298606
rect 187263 298578 187291 298606
rect 187077 298516 187105 298544
rect 187139 298516 187167 298544
rect 187201 298516 187229 298544
rect 187263 298516 187291 298544
rect 187077 298454 187105 298482
rect 187139 298454 187167 298482
rect 187201 298454 187229 298482
rect 187263 298454 187291 298482
rect 187077 298392 187105 298420
rect 187139 298392 187167 298420
rect 187201 298392 187229 298420
rect 187263 298392 187291 298420
rect 187077 290147 187105 290175
rect 187139 290147 187167 290175
rect 187201 290147 187229 290175
rect 187263 290147 187291 290175
rect 187077 290085 187105 290113
rect 187139 290085 187167 290113
rect 187201 290085 187229 290113
rect 187263 290085 187291 290113
rect 187077 290023 187105 290051
rect 187139 290023 187167 290051
rect 187201 290023 187229 290051
rect 187263 290023 187291 290051
rect 187077 289961 187105 289989
rect 187139 289961 187167 289989
rect 187201 289961 187229 289989
rect 187263 289961 187291 289989
rect 187077 281147 187105 281175
rect 187139 281147 187167 281175
rect 187201 281147 187229 281175
rect 187263 281147 187291 281175
rect 187077 281085 187105 281113
rect 187139 281085 187167 281113
rect 187201 281085 187229 281113
rect 187263 281085 187291 281113
rect 187077 281023 187105 281051
rect 187139 281023 187167 281051
rect 187201 281023 187229 281051
rect 187263 281023 187291 281051
rect 187077 280961 187105 280989
rect 187139 280961 187167 280989
rect 187201 280961 187229 280989
rect 187263 280961 187291 280989
rect 187077 272147 187105 272175
rect 187139 272147 187167 272175
rect 187201 272147 187229 272175
rect 187263 272147 187291 272175
rect 187077 272085 187105 272113
rect 187139 272085 187167 272113
rect 187201 272085 187229 272113
rect 187263 272085 187291 272113
rect 187077 272023 187105 272051
rect 187139 272023 187167 272051
rect 187201 272023 187229 272051
rect 187263 272023 187291 272051
rect 187077 271961 187105 271989
rect 187139 271961 187167 271989
rect 187201 271961 187229 271989
rect 187263 271961 187291 271989
rect 187077 263147 187105 263175
rect 187139 263147 187167 263175
rect 187201 263147 187229 263175
rect 187263 263147 187291 263175
rect 187077 263085 187105 263113
rect 187139 263085 187167 263113
rect 187201 263085 187229 263113
rect 187263 263085 187291 263113
rect 187077 263023 187105 263051
rect 187139 263023 187167 263051
rect 187201 263023 187229 263051
rect 187263 263023 187291 263051
rect 187077 262961 187105 262989
rect 187139 262961 187167 262989
rect 187201 262961 187229 262989
rect 187263 262961 187291 262989
rect 187077 254147 187105 254175
rect 187139 254147 187167 254175
rect 187201 254147 187229 254175
rect 187263 254147 187291 254175
rect 187077 254085 187105 254113
rect 187139 254085 187167 254113
rect 187201 254085 187229 254113
rect 187263 254085 187291 254113
rect 187077 254023 187105 254051
rect 187139 254023 187167 254051
rect 187201 254023 187229 254051
rect 187263 254023 187291 254051
rect 187077 253961 187105 253989
rect 187139 253961 187167 253989
rect 187201 253961 187229 253989
rect 187263 253961 187291 253989
rect 187077 245147 187105 245175
rect 187139 245147 187167 245175
rect 187201 245147 187229 245175
rect 187263 245147 187291 245175
rect 187077 245085 187105 245113
rect 187139 245085 187167 245113
rect 187201 245085 187229 245113
rect 187263 245085 187291 245113
rect 187077 245023 187105 245051
rect 187139 245023 187167 245051
rect 187201 245023 187229 245051
rect 187263 245023 187291 245051
rect 187077 244961 187105 244989
rect 187139 244961 187167 244989
rect 187201 244961 187229 244989
rect 187263 244961 187291 244989
rect 187077 236147 187105 236175
rect 187139 236147 187167 236175
rect 187201 236147 187229 236175
rect 187263 236147 187291 236175
rect 187077 236085 187105 236113
rect 187139 236085 187167 236113
rect 187201 236085 187229 236113
rect 187263 236085 187291 236113
rect 187077 236023 187105 236051
rect 187139 236023 187167 236051
rect 187201 236023 187229 236051
rect 187263 236023 187291 236051
rect 187077 235961 187105 235989
rect 187139 235961 187167 235989
rect 187201 235961 187229 235989
rect 187263 235961 187291 235989
rect 187077 227147 187105 227175
rect 187139 227147 187167 227175
rect 187201 227147 187229 227175
rect 187263 227147 187291 227175
rect 187077 227085 187105 227113
rect 187139 227085 187167 227113
rect 187201 227085 187229 227113
rect 187263 227085 187291 227113
rect 187077 227023 187105 227051
rect 187139 227023 187167 227051
rect 187201 227023 187229 227051
rect 187263 227023 187291 227051
rect 187077 226961 187105 226989
rect 187139 226961 187167 226989
rect 187201 226961 187229 226989
rect 187263 226961 187291 226989
rect 187077 218147 187105 218175
rect 187139 218147 187167 218175
rect 187201 218147 187229 218175
rect 187263 218147 187291 218175
rect 187077 218085 187105 218113
rect 187139 218085 187167 218113
rect 187201 218085 187229 218113
rect 187263 218085 187291 218113
rect 187077 218023 187105 218051
rect 187139 218023 187167 218051
rect 187201 218023 187229 218051
rect 187263 218023 187291 218051
rect 187077 217961 187105 217989
rect 187139 217961 187167 217989
rect 187201 217961 187229 217989
rect 187263 217961 187291 217989
rect 187077 209147 187105 209175
rect 187139 209147 187167 209175
rect 187201 209147 187229 209175
rect 187263 209147 187291 209175
rect 187077 209085 187105 209113
rect 187139 209085 187167 209113
rect 187201 209085 187229 209113
rect 187263 209085 187291 209113
rect 187077 209023 187105 209051
rect 187139 209023 187167 209051
rect 187201 209023 187229 209051
rect 187263 209023 187291 209051
rect 187077 208961 187105 208989
rect 187139 208961 187167 208989
rect 187201 208961 187229 208989
rect 187263 208961 187291 208989
rect 187077 200147 187105 200175
rect 187139 200147 187167 200175
rect 187201 200147 187229 200175
rect 187263 200147 187291 200175
rect 187077 200085 187105 200113
rect 187139 200085 187167 200113
rect 187201 200085 187229 200113
rect 187263 200085 187291 200113
rect 187077 200023 187105 200051
rect 187139 200023 187167 200051
rect 187201 200023 187229 200051
rect 187263 200023 187291 200051
rect 187077 199961 187105 199989
rect 187139 199961 187167 199989
rect 187201 199961 187229 199989
rect 187263 199961 187291 199989
rect 188937 299058 188965 299086
rect 188999 299058 189027 299086
rect 189061 299058 189089 299086
rect 189123 299058 189151 299086
rect 188937 298996 188965 299024
rect 188999 298996 189027 299024
rect 189061 298996 189089 299024
rect 189123 298996 189151 299024
rect 188937 298934 188965 298962
rect 188999 298934 189027 298962
rect 189061 298934 189089 298962
rect 189123 298934 189151 298962
rect 188937 298872 188965 298900
rect 188999 298872 189027 298900
rect 189061 298872 189089 298900
rect 189123 298872 189151 298900
rect 188937 293147 188965 293175
rect 188999 293147 189027 293175
rect 189061 293147 189089 293175
rect 189123 293147 189151 293175
rect 188937 293085 188965 293113
rect 188999 293085 189027 293113
rect 189061 293085 189089 293113
rect 189123 293085 189151 293113
rect 188937 293023 188965 293051
rect 188999 293023 189027 293051
rect 189061 293023 189089 293051
rect 189123 293023 189151 293051
rect 188937 292961 188965 292989
rect 188999 292961 189027 292989
rect 189061 292961 189089 292989
rect 189123 292961 189151 292989
rect 188937 284147 188965 284175
rect 188999 284147 189027 284175
rect 189061 284147 189089 284175
rect 189123 284147 189151 284175
rect 188937 284085 188965 284113
rect 188999 284085 189027 284113
rect 189061 284085 189089 284113
rect 189123 284085 189151 284113
rect 188937 284023 188965 284051
rect 188999 284023 189027 284051
rect 189061 284023 189089 284051
rect 189123 284023 189151 284051
rect 188937 283961 188965 283989
rect 188999 283961 189027 283989
rect 189061 283961 189089 283989
rect 189123 283961 189151 283989
rect 188937 275147 188965 275175
rect 188999 275147 189027 275175
rect 189061 275147 189089 275175
rect 189123 275147 189151 275175
rect 188937 275085 188965 275113
rect 188999 275085 189027 275113
rect 189061 275085 189089 275113
rect 189123 275085 189151 275113
rect 188937 275023 188965 275051
rect 188999 275023 189027 275051
rect 189061 275023 189089 275051
rect 189123 275023 189151 275051
rect 188937 274961 188965 274989
rect 188999 274961 189027 274989
rect 189061 274961 189089 274989
rect 189123 274961 189151 274989
rect 188937 266147 188965 266175
rect 188999 266147 189027 266175
rect 189061 266147 189089 266175
rect 189123 266147 189151 266175
rect 188937 266085 188965 266113
rect 188999 266085 189027 266113
rect 189061 266085 189089 266113
rect 189123 266085 189151 266113
rect 188937 266023 188965 266051
rect 188999 266023 189027 266051
rect 189061 266023 189089 266051
rect 189123 266023 189151 266051
rect 188937 265961 188965 265989
rect 188999 265961 189027 265989
rect 189061 265961 189089 265989
rect 189123 265961 189151 265989
rect 188937 257147 188965 257175
rect 188999 257147 189027 257175
rect 189061 257147 189089 257175
rect 189123 257147 189151 257175
rect 188937 257085 188965 257113
rect 188999 257085 189027 257113
rect 189061 257085 189089 257113
rect 189123 257085 189151 257113
rect 188937 257023 188965 257051
rect 188999 257023 189027 257051
rect 189061 257023 189089 257051
rect 189123 257023 189151 257051
rect 188937 256961 188965 256989
rect 188999 256961 189027 256989
rect 189061 256961 189089 256989
rect 189123 256961 189151 256989
rect 188937 248147 188965 248175
rect 188999 248147 189027 248175
rect 189061 248147 189089 248175
rect 189123 248147 189151 248175
rect 188937 248085 188965 248113
rect 188999 248085 189027 248113
rect 189061 248085 189089 248113
rect 189123 248085 189151 248113
rect 188937 248023 188965 248051
rect 188999 248023 189027 248051
rect 189061 248023 189089 248051
rect 189123 248023 189151 248051
rect 188937 247961 188965 247989
rect 188999 247961 189027 247989
rect 189061 247961 189089 247989
rect 189123 247961 189151 247989
rect 188937 239147 188965 239175
rect 188999 239147 189027 239175
rect 189061 239147 189089 239175
rect 189123 239147 189151 239175
rect 188937 239085 188965 239113
rect 188999 239085 189027 239113
rect 189061 239085 189089 239113
rect 189123 239085 189151 239113
rect 188937 239023 188965 239051
rect 188999 239023 189027 239051
rect 189061 239023 189089 239051
rect 189123 239023 189151 239051
rect 188937 238961 188965 238989
rect 188999 238961 189027 238989
rect 189061 238961 189089 238989
rect 189123 238961 189151 238989
rect 188937 230147 188965 230175
rect 188999 230147 189027 230175
rect 189061 230147 189089 230175
rect 189123 230147 189151 230175
rect 188937 230085 188965 230113
rect 188999 230085 189027 230113
rect 189061 230085 189089 230113
rect 189123 230085 189151 230113
rect 188937 230023 188965 230051
rect 188999 230023 189027 230051
rect 189061 230023 189089 230051
rect 189123 230023 189151 230051
rect 188937 229961 188965 229989
rect 188999 229961 189027 229989
rect 189061 229961 189089 229989
rect 189123 229961 189151 229989
rect 188937 221147 188965 221175
rect 188999 221147 189027 221175
rect 189061 221147 189089 221175
rect 189123 221147 189151 221175
rect 188937 221085 188965 221113
rect 188999 221085 189027 221113
rect 189061 221085 189089 221113
rect 189123 221085 189151 221113
rect 188937 221023 188965 221051
rect 188999 221023 189027 221051
rect 189061 221023 189089 221051
rect 189123 221023 189151 221051
rect 188937 220961 188965 220989
rect 188999 220961 189027 220989
rect 189061 220961 189089 220989
rect 189123 220961 189151 220989
rect 188937 212147 188965 212175
rect 188999 212147 189027 212175
rect 189061 212147 189089 212175
rect 189123 212147 189151 212175
rect 188937 212085 188965 212113
rect 188999 212085 189027 212113
rect 189061 212085 189089 212113
rect 189123 212085 189151 212113
rect 188937 212023 188965 212051
rect 188999 212023 189027 212051
rect 189061 212023 189089 212051
rect 189123 212023 189151 212051
rect 188937 211961 188965 211989
rect 188999 211961 189027 211989
rect 189061 211961 189089 211989
rect 189123 211961 189151 211989
rect 188937 203147 188965 203175
rect 188999 203147 189027 203175
rect 189061 203147 189089 203175
rect 189123 203147 189151 203175
rect 188937 203085 188965 203113
rect 188999 203085 189027 203113
rect 189061 203085 189089 203113
rect 189123 203085 189151 203113
rect 188937 203023 188965 203051
rect 188999 203023 189027 203051
rect 189061 203023 189089 203051
rect 189123 203023 189151 203051
rect 188937 202961 188965 202989
rect 188999 202961 189027 202989
rect 189061 202961 189089 202989
rect 189123 202961 189151 202989
rect 202437 298578 202465 298606
rect 202499 298578 202527 298606
rect 202561 298578 202589 298606
rect 202623 298578 202651 298606
rect 202437 298516 202465 298544
rect 202499 298516 202527 298544
rect 202561 298516 202589 298544
rect 202623 298516 202651 298544
rect 202437 298454 202465 298482
rect 202499 298454 202527 298482
rect 202561 298454 202589 298482
rect 202623 298454 202651 298482
rect 202437 298392 202465 298420
rect 202499 298392 202527 298420
rect 202561 298392 202589 298420
rect 202623 298392 202651 298420
rect 202437 290147 202465 290175
rect 202499 290147 202527 290175
rect 202561 290147 202589 290175
rect 202623 290147 202651 290175
rect 202437 290085 202465 290113
rect 202499 290085 202527 290113
rect 202561 290085 202589 290113
rect 202623 290085 202651 290113
rect 202437 290023 202465 290051
rect 202499 290023 202527 290051
rect 202561 290023 202589 290051
rect 202623 290023 202651 290051
rect 202437 289961 202465 289989
rect 202499 289961 202527 289989
rect 202561 289961 202589 289989
rect 202623 289961 202651 289989
rect 202437 281147 202465 281175
rect 202499 281147 202527 281175
rect 202561 281147 202589 281175
rect 202623 281147 202651 281175
rect 202437 281085 202465 281113
rect 202499 281085 202527 281113
rect 202561 281085 202589 281113
rect 202623 281085 202651 281113
rect 202437 281023 202465 281051
rect 202499 281023 202527 281051
rect 202561 281023 202589 281051
rect 202623 281023 202651 281051
rect 202437 280961 202465 280989
rect 202499 280961 202527 280989
rect 202561 280961 202589 280989
rect 202623 280961 202651 280989
rect 202437 272147 202465 272175
rect 202499 272147 202527 272175
rect 202561 272147 202589 272175
rect 202623 272147 202651 272175
rect 202437 272085 202465 272113
rect 202499 272085 202527 272113
rect 202561 272085 202589 272113
rect 202623 272085 202651 272113
rect 202437 272023 202465 272051
rect 202499 272023 202527 272051
rect 202561 272023 202589 272051
rect 202623 272023 202651 272051
rect 202437 271961 202465 271989
rect 202499 271961 202527 271989
rect 202561 271961 202589 271989
rect 202623 271961 202651 271989
rect 202437 263147 202465 263175
rect 202499 263147 202527 263175
rect 202561 263147 202589 263175
rect 202623 263147 202651 263175
rect 202437 263085 202465 263113
rect 202499 263085 202527 263113
rect 202561 263085 202589 263113
rect 202623 263085 202651 263113
rect 202437 263023 202465 263051
rect 202499 263023 202527 263051
rect 202561 263023 202589 263051
rect 202623 263023 202651 263051
rect 202437 262961 202465 262989
rect 202499 262961 202527 262989
rect 202561 262961 202589 262989
rect 202623 262961 202651 262989
rect 202437 254147 202465 254175
rect 202499 254147 202527 254175
rect 202561 254147 202589 254175
rect 202623 254147 202651 254175
rect 202437 254085 202465 254113
rect 202499 254085 202527 254113
rect 202561 254085 202589 254113
rect 202623 254085 202651 254113
rect 202437 254023 202465 254051
rect 202499 254023 202527 254051
rect 202561 254023 202589 254051
rect 202623 254023 202651 254051
rect 202437 253961 202465 253989
rect 202499 253961 202527 253989
rect 202561 253961 202589 253989
rect 202623 253961 202651 253989
rect 202437 245147 202465 245175
rect 202499 245147 202527 245175
rect 202561 245147 202589 245175
rect 202623 245147 202651 245175
rect 202437 245085 202465 245113
rect 202499 245085 202527 245113
rect 202561 245085 202589 245113
rect 202623 245085 202651 245113
rect 202437 245023 202465 245051
rect 202499 245023 202527 245051
rect 202561 245023 202589 245051
rect 202623 245023 202651 245051
rect 202437 244961 202465 244989
rect 202499 244961 202527 244989
rect 202561 244961 202589 244989
rect 202623 244961 202651 244989
rect 202437 236147 202465 236175
rect 202499 236147 202527 236175
rect 202561 236147 202589 236175
rect 202623 236147 202651 236175
rect 202437 236085 202465 236113
rect 202499 236085 202527 236113
rect 202561 236085 202589 236113
rect 202623 236085 202651 236113
rect 202437 236023 202465 236051
rect 202499 236023 202527 236051
rect 202561 236023 202589 236051
rect 202623 236023 202651 236051
rect 202437 235961 202465 235989
rect 202499 235961 202527 235989
rect 202561 235961 202589 235989
rect 202623 235961 202651 235989
rect 202437 227147 202465 227175
rect 202499 227147 202527 227175
rect 202561 227147 202589 227175
rect 202623 227147 202651 227175
rect 202437 227085 202465 227113
rect 202499 227085 202527 227113
rect 202561 227085 202589 227113
rect 202623 227085 202651 227113
rect 202437 227023 202465 227051
rect 202499 227023 202527 227051
rect 202561 227023 202589 227051
rect 202623 227023 202651 227051
rect 202437 226961 202465 226989
rect 202499 226961 202527 226989
rect 202561 226961 202589 226989
rect 202623 226961 202651 226989
rect 202437 218147 202465 218175
rect 202499 218147 202527 218175
rect 202561 218147 202589 218175
rect 202623 218147 202651 218175
rect 202437 218085 202465 218113
rect 202499 218085 202527 218113
rect 202561 218085 202589 218113
rect 202623 218085 202651 218113
rect 202437 218023 202465 218051
rect 202499 218023 202527 218051
rect 202561 218023 202589 218051
rect 202623 218023 202651 218051
rect 202437 217961 202465 217989
rect 202499 217961 202527 217989
rect 202561 217961 202589 217989
rect 202623 217961 202651 217989
rect 202437 209147 202465 209175
rect 202499 209147 202527 209175
rect 202561 209147 202589 209175
rect 202623 209147 202651 209175
rect 202437 209085 202465 209113
rect 202499 209085 202527 209113
rect 202561 209085 202589 209113
rect 202623 209085 202651 209113
rect 202437 209023 202465 209051
rect 202499 209023 202527 209051
rect 202561 209023 202589 209051
rect 202623 209023 202651 209051
rect 202437 208961 202465 208989
rect 202499 208961 202527 208989
rect 202561 208961 202589 208989
rect 202623 208961 202651 208989
rect 202437 200147 202465 200175
rect 202499 200147 202527 200175
rect 202561 200147 202589 200175
rect 202623 200147 202651 200175
rect 202437 200085 202465 200113
rect 202499 200085 202527 200113
rect 202561 200085 202589 200113
rect 202623 200085 202651 200113
rect 202437 200023 202465 200051
rect 202499 200023 202527 200051
rect 202561 200023 202589 200051
rect 202623 200023 202651 200051
rect 202437 199961 202465 199989
rect 202499 199961 202527 199989
rect 202561 199961 202589 199989
rect 202623 199961 202651 199989
rect 188937 194147 188965 194175
rect 188999 194147 189027 194175
rect 189061 194147 189089 194175
rect 189123 194147 189151 194175
rect 188937 194085 188965 194113
rect 188999 194085 189027 194113
rect 189061 194085 189089 194113
rect 189123 194085 189151 194113
rect 188937 194023 188965 194051
rect 188999 194023 189027 194051
rect 189061 194023 189089 194051
rect 189123 194023 189151 194051
rect 188937 193961 188965 193989
rect 188999 193961 189027 193989
rect 189061 193961 189089 193989
rect 189123 193961 189151 193989
rect 189939 194147 189967 194175
rect 190001 194147 190029 194175
rect 189939 194085 189967 194113
rect 190001 194085 190029 194113
rect 189939 194023 189967 194051
rect 190001 194023 190029 194051
rect 189939 193961 189967 193989
rect 190001 193961 190029 193989
rect 182259 191147 182287 191175
rect 182321 191147 182349 191175
rect 182259 191085 182287 191113
rect 182321 191085 182349 191113
rect 182259 191023 182287 191051
rect 182321 191023 182349 191051
rect 182259 190961 182287 190989
rect 182321 190961 182349 190989
rect 197619 191147 197647 191175
rect 197681 191147 197709 191175
rect 197619 191085 197647 191113
rect 197681 191085 197709 191113
rect 197619 191023 197647 191051
rect 197681 191023 197709 191051
rect 197619 190961 197647 190989
rect 197681 190961 197709 190989
rect 202437 191147 202465 191175
rect 202499 191147 202527 191175
rect 202561 191147 202589 191175
rect 202623 191147 202651 191175
rect 202437 191085 202465 191113
rect 202499 191085 202527 191113
rect 202561 191085 202589 191113
rect 202623 191085 202651 191113
rect 202437 191023 202465 191051
rect 202499 191023 202527 191051
rect 202561 191023 202589 191051
rect 202623 191023 202651 191051
rect 202437 190961 202465 190989
rect 202499 190961 202527 190989
rect 202561 190961 202589 190989
rect 202623 190961 202651 190989
rect 173577 185147 173605 185175
rect 173639 185147 173667 185175
rect 173701 185147 173729 185175
rect 173763 185147 173791 185175
rect 173577 185085 173605 185113
rect 173639 185085 173667 185113
rect 173701 185085 173729 185113
rect 173763 185085 173791 185113
rect 173577 185023 173605 185051
rect 173639 185023 173667 185051
rect 173701 185023 173729 185051
rect 173763 185023 173791 185051
rect 173577 184961 173605 184989
rect 173639 184961 173667 184989
rect 173701 184961 173729 184989
rect 173763 184961 173791 184989
rect 189939 185147 189967 185175
rect 190001 185147 190029 185175
rect 189939 185085 189967 185113
rect 190001 185085 190029 185113
rect 189939 185023 189967 185051
rect 190001 185023 190029 185051
rect 189939 184961 189967 184989
rect 190001 184961 190029 184989
rect 182259 182147 182287 182175
rect 182321 182147 182349 182175
rect 182259 182085 182287 182113
rect 182321 182085 182349 182113
rect 182259 182023 182287 182051
rect 182321 182023 182349 182051
rect 182259 181961 182287 181989
rect 182321 181961 182349 181989
rect 197619 182147 197647 182175
rect 197681 182147 197709 182175
rect 197619 182085 197647 182113
rect 197681 182085 197709 182113
rect 197619 182023 197647 182051
rect 197681 182023 197709 182051
rect 197619 181961 197647 181989
rect 197681 181961 197709 181989
rect 202437 182147 202465 182175
rect 202499 182147 202527 182175
rect 202561 182147 202589 182175
rect 202623 182147 202651 182175
rect 202437 182085 202465 182113
rect 202499 182085 202527 182113
rect 202561 182085 202589 182113
rect 202623 182085 202651 182113
rect 202437 182023 202465 182051
rect 202499 182023 202527 182051
rect 202561 182023 202589 182051
rect 202623 182023 202651 182051
rect 202437 181961 202465 181989
rect 202499 181961 202527 181989
rect 202561 181961 202589 181989
rect 202623 181961 202651 181989
rect 173577 176147 173605 176175
rect 173639 176147 173667 176175
rect 173701 176147 173729 176175
rect 173763 176147 173791 176175
rect 173577 176085 173605 176113
rect 173639 176085 173667 176113
rect 173701 176085 173729 176113
rect 173763 176085 173791 176113
rect 173577 176023 173605 176051
rect 173639 176023 173667 176051
rect 173701 176023 173729 176051
rect 173763 176023 173791 176051
rect 173577 175961 173605 175989
rect 173639 175961 173667 175989
rect 173701 175961 173729 175989
rect 173763 175961 173791 175989
rect 189939 176147 189967 176175
rect 190001 176147 190029 176175
rect 189939 176085 189967 176113
rect 190001 176085 190029 176113
rect 189939 176023 189967 176051
rect 190001 176023 190029 176051
rect 189939 175961 189967 175989
rect 190001 175961 190029 175989
rect 182259 173147 182287 173175
rect 182321 173147 182349 173175
rect 182259 173085 182287 173113
rect 182321 173085 182349 173113
rect 182259 173023 182287 173051
rect 182321 173023 182349 173051
rect 182259 172961 182287 172989
rect 182321 172961 182349 172989
rect 187077 173147 187105 173175
rect 187139 173147 187167 173175
rect 187201 173147 187229 173175
rect 187263 173147 187291 173175
rect 187077 173085 187105 173113
rect 187139 173085 187167 173113
rect 187201 173085 187229 173113
rect 187263 173085 187291 173113
rect 187077 173023 187105 173051
rect 187139 173023 187167 173051
rect 187201 173023 187229 173051
rect 187263 173023 187291 173051
rect 187077 172961 187105 172989
rect 187139 172961 187167 172989
rect 187201 172961 187229 172989
rect 187263 172961 187291 172989
rect 173577 167147 173605 167175
rect 173639 167147 173667 167175
rect 173701 167147 173729 167175
rect 173763 167147 173791 167175
rect 173577 167085 173605 167113
rect 173639 167085 173667 167113
rect 173701 167085 173729 167113
rect 173763 167085 173791 167113
rect 173577 167023 173605 167051
rect 173639 167023 173667 167051
rect 173701 167023 173729 167051
rect 173763 167023 173791 167051
rect 173577 166961 173605 166989
rect 173639 166961 173667 166989
rect 173701 166961 173729 166989
rect 173763 166961 173791 166989
rect 197619 173147 197647 173175
rect 197681 173147 197709 173175
rect 197619 173085 197647 173113
rect 197681 173085 197709 173113
rect 197619 173023 197647 173051
rect 197681 173023 197709 173051
rect 197619 172961 197647 172989
rect 197681 172961 197709 172989
rect 202437 173147 202465 173175
rect 202499 173147 202527 173175
rect 202561 173147 202589 173175
rect 202623 173147 202651 173175
rect 202437 173085 202465 173113
rect 202499 173085 202527 173113
rect 202561 173085 202589 173113
rect 202623 173085 202651 173113
rect 202437 173023 202465 173051
rect 202499 173023 202527 173051
rect 202561 173023 202589 173051
rect 202623 173023 202651 173051
rect 202437 172961 202465 172989
rect 202499 172961 202527 172989
rect 202561 172961 202589 172989
rect 202623 172961 202651 172989
rect 187077 164147 187105 164175
rect 187139 164147 187167 164175
rect 187201 164147 187229 164175
rect 187263 164147 187291 164175
rect 187077 164085 187105 164113
rect 187139 164085 187167 164113
rect 187201 164085 187229 164113
rect 187263 164085 187291 164113
rect 187077 164023 187105 164051
rect 187139 164023 187167 164051
rect 187201 164023 187229 164051
rect 187263 164023 187291 164051
rect 187077 163961 187105 163989
rect 187139 163961 187167 163989
rect 187201 163961 187229 163989
rect 187263 163961 187291 163989
rect 202437 164147 202465 164175
rect 202499 164147 202527 164175
rect 202561 164147 202589 164175
rect 202623 164147 202651 164175
rect 202437 164085 202465 164113
rect 202499 164085 202527 164113
rect 202561 164085 202589 164113
rect 202623 164085 202651 164113
rect 202437 164023 202465 164051
rect 202499 164023 202527 164051
rect 202561 164023 202589 164051
rect 202623 164023 202651 164051
rect 202437 163961 202465 163989
rect 202499 163961 202527 163989
rect 202561 163961 202589 163989
rect 202623 163961 202651 163989
rect 204297 299058 204325 299086
rect 204359 299058 204387 299086
rect 204421 299058 204449 299086
rect 204483 299058 204511 299086
rect 204297 298996 204325 299024
rect 204359 298996 204387 299024
rect 204421 298996 204449 299024
rect 204483 298996 204511 299024
rect 204297 298934 204325 298962
rect 204359 298934 204387 298962
rect 204421 298934 204449 298962
rect 204483 298934 204511 298962
rect 204297 298872 204325 298900
rect 204359 298872 204387 298900
rect 204421 298872 204449 298900
rect 204483 298872 204511 298900
rect 204297 293147 204325 293175
rect 204359 293147 204387 293175
rect 204421 293147 204449 293175
rect 204483 293147 204511 293175
rect 204297 293085 204325 293113
rect 204359 293085 204387 293113
rect 204421 293085 204449 293113
rect 204483 293085 204511 293113
rect 204297 293023 204325 293051
rect 204359 293023 204387 293051
rect 204421 293023 204449 293051
rect 204483 293023 204511 293051
rect 204297 292961 204325 292989
rect 204359 292961 204387 292989
rect 204421 292961 204449 292989
rect 204483 292961 204511 292989
rect 204297 284147 204325 284175
rect 204359 284147 204387 284175
rect 204421 284147 204449 284175
rect 204483 284147 204511 284175
rect 204297 284085 204325 284113
rect 204359 284085 204387 284113
rect 204421 284085 204449 284113
rect 204483 284085 204511 284113
rect 204297 284023 204325 284051
rect 204359 284023 204387 284051
rect 204421 284023 204449 284051
rect 204483 284023 204511 284051
rect 204297 283961 204325 283989
rect 204359 283961 204387 283989
rect 204421 283961 204449 283989
rect 204483 283961 204511 283989
rect 204297 275147 204325 275175
rect 204359 275147 204387 275175
rect 204421 275147 204449 275175
rect 204483 275147 204511 275175
rect 204297 275085 204325 275113
rect 204359 275085 204387 275113
rect 204421 275085 204449 275113
rect 204483 275085 204511 275113
rect 204297 275023 204325 275051
rect 204359 275023 204387 275051
rect 204421 275023 204449 275051
rect 204483 275023 204511 275051
rect 204297 274961 204325 274989
rect 204359 274961 204387 274989
rect 204421 274961 204449 274989
rect 204483 274961 204511 274989
rect 204297 266147 204325 266175
rect 204359 266147 204387 266175
rect 204421 266147 204449 266175
rect 204483 266147 204511 266175
rect 204297 266085 204325 266113
rect 204359 266085 204387 266113
rect 204421 266085 204449 266113
rect 204483 266085 204511 266113
rect 204297 266023 204325 266051
rect 204359 266023 204387 266051
rect 204421 266023 204449 266051
rect 204483 266023 204511 266051
rect 204297 265961 204325 265989
rect 204359 265961 204387 265989
rect 204421 265961 204449 265989
rect 204483 265961 204511 265989
rect 204297 257147 204325 257175
rect 204359 257147 204387 257175
rect 204421 257147 204449 257175
rect 204483 257147 204511 257175
rect 204297 257085 204325 257113
rect 204359 257085 204387 257113
rect 204421 257085 204449 257113
rect 204483 257085 204511 257113
rect 204297 257023 204325 257051
rect 204359 257023 204387 257051
rect 204421 257023 204449 257051
rect 204483 257023 204511 257051
rect 204297 256961 204325 256989
rect 204359 256961 204387 256989
rect 204421 256961 204449 256989
rect 204483 256961 204511 256989
rect 204297 248147 204325 248175
rect 204359 248147 204387 248175
rect 204421 248147 204449 248175
rect 204483 248147 204511 248175
rect 204297 248085 204325 248113
rect 204359 248085 204387 248113
rect 204421 248085 204449 248113
rect 204483 248085 204511 248113
rect 204297 248023 204325 248051
rect 204359 248023 204387 248051
rect 204421 248023 204449 248051
rect 204483 248023 204511 248051
rect 204297 247961 204325 247989
rect 204359 247961 204387 247989
rect 204421 247961 204449 247989
rect 204483 247961 204511 247989
rect 204297 239147 204325 239175
rect 204359 239147 204387 239175
rect 204421 239147 204449 239175
rect 204483 239147 204511 239175
rect 204297 239085 204325 239113
rect 204359 239085 204387 239113
rect 204421 239085 204449 239113
rect 204483 239085 204511 239113
rect 204297 239023 204325 239051
rect 204359 239023 204387 239051
rect 204421 239023 204449 239051
rect 204483 239023 204511 239051
rect 204297 238961 204325 238989
rect 204359 238961 204387 238989
rect 204421 238961 204449 238989
rect 204483 238961 204511 238989
rect 204297 230147 204325 230175
rect 204359 230147 204387 230175
rect 204421 230147 204449 230175
rect 204483 230147 204511 230175
rect 204297 230085 204325 230113
rect 204359 230085 204387 230113
rect 204421 230085 204449 230113
rect 204483 230085 204511 230113
rect 204297 230023 204325 230051
rect 204359 230023 204387 230051
rect 204421 230023 204449 230051
rect 204483 230023 204511 230051
rect 204297 229961 204325 229989
rect 204359 229961 204387 229989
rect 204421 229961 204449 229989
rect 204483 229961 204511 229989
rect 204297 221147 204325 221175
rect 204359 221147 204387 221175
rect 204421 221147 204449 221175
rect 204483 221147 204511 221175
rect 204297 221085 204325 221113
rect 204359 221085 204387 221113
rect 204421 221085 204449 221113
rect 204483 221085 204511 221113
rect 204297 221023 204325 221051
rect 204359 221023 204387 221051
rect 204421 221023 204449 221051
rect 204483 221023 204511 221051
rect 204297 220961 204325 220989
rect 204359 220961 204387 220989
rect 204421 220961 204449 220989
rect 204483 220961 204511 220989
rect 204297 212147 204325 212175
rect 204359 212147 204387 212175
rect 204421 212147 204449 212175
rect 204483 212147 204511 212175
rect 204297 212085 204325 212113
rect 204359 212085 204387 212113
rect 204421 212085 204449 212113
rect 204483 212085 204511 212113
rect 204297 212023 204325 212051
rect 204359 212023 204387 212051
rect 204421 212023 204449 212051
rect 204483 212023 204511 212051
rect 204297 211961 204325 211989
rect 204359 211961 204387 211989
rect 204421 211961 204449 211989
rect 204483 211961 204511 211989
rect 204297 203147 204325 203175
rect 204359 203147 204387 203175
rect 204421 203147 204449 203175
rect 204483 203147 204511 203175
rect 204297 203085 204325 203113
rect 204359 203085 204387 203113
rect 204421 203085 204449 203113
rect 204483 203085 204511 203113
rect 204297 203023 204325 203051
rect 204359 203023 204387 203051
rect 204421 203023 204449 203051
rect 204483 203023 204511 203051
rect 204297 202961 204325 202989
rect 204359 202961 204387 202989
rect 204421 202961 204449 202989
rect 204483 202961 204511 202989
rect 204297 194147 204325 194175
rect 204359 194147 204387 194175
rect 204421 194147 204449 194175
rect 204483 194147 204511 194175
rect 204297 194085 204325 194113
rect 204359 194085 204387 194113
rect 204421 194085 204449 194113
rect 204483 194085 204511 194113
rect 204297 194023 204325 194051
rect 204359 194023 204387 194051
rect 204421 194023 204449 194051
rect 204483 194023 204511 194051
rect 204297 193961 204325 193989
rect 204359 193961 204387 193989
rect 204421 193961 204449 193989
rect 204483 193961 204511 193989
rect 204297 185147 204325 185175
rect 204359 185147 204387 185175
rect 204421 185147 204449 185175
rect 204483 185147 204511 185175
rect 204297 185085 204325 185113
rect 204359 185085 204387 185113
rect 204421 185085 204449 185113
rect 204483 185085 204511 185113
rect 204297 185023 204325 185051
rect 204359 185023 204387 185051
rect 204421 185023 204449 185051
rect 204483 185023 204511 185051
rect 204297 184961 204325 184989
rect 204359 184961 204387 184989
rect 204421 184961 204449 184989
rect 204483 184961 204511 184989
rect 204297 176147 204325 176175
rect 204359 176147 204387 176175
rect 204421 176147 204449 176175
rect 204483 176147 204511 176175
rect 204297 176085 204325 176113
rect 204359 176085 204387 176113
rect 204421 176085 204449 176113
rect 204483 176085 204511 176113
rect 204297 176023 204325 176051
rect 204359 176023 204387 176051
rect 204421 176023 204449 176051
rect 204483 176023 204511 176051
rect 204297 175961 204325 175989
rect 204359 175961 204387 175989
rect 204421 175961 204449 175989
rect 204483 175961 204511 175989
rect 204297 167147 204325 167175
rect 204359 167147 204387 167175
rect 204421 167147 204449 167175
rect 204483 167147 204511 167175
rect 204297 167085 204325 167113
rect 204359 167085 204387 167113
rect 204421 167085 204449 167113
rect 204483 167085 204511 167113
rect 204297 167023 204325 167051
rect 204359 167023 204387 167051
rect 204421 167023 204449 167051
rect 204483 167023 204511 167051
rect 204297 166961 204325 166989
rect 204359 166961 204387 166989
rect 204421 166961 204449 166989
rect 204483 166961 204511 166989
rect 96777 158147 96805 158175
rect 96839 158147 96867 158175
rect 96901 158147 96929 158175
rect 96963 158147 96991 158175
rect 96777 158085 96805 158113
rect 96839 158085 96867 158113
rect 96901 158085 96929 158113
rect 96963 158085 96991 158113
rect 96777 158023 96805 158051
rect 96839 158023 96867 158051
rect 96901 158023 96929 158051
rect 96963 158023 96991 158051
rect 96777 157961 96805 157989
rect 96839 157961 96867 157989
rect 96901 157961 96929 157989
rect 96963 157961 96991 157989
rect 101379 158147 101407 158175
rect 101441 158147 101469 158175
rect 101379 158085 101407 158113
rect 101441 158085 101469 158113
rect 101379 158023 101407 158051
rect 101441 158023 101469 158051
rect 101379 157961 101407 157989
rect 101441 157961 101469 157989
rect 116739 158147 116767 158175
rect 116801 158147 116829 158175
rect 116739 158085 116767 158113
rect 116801 158085 116829 158113
rect 116739 158023 116767 158051
rect 116801 158023 116829 158051
rect 116739 157961 116767 157989
rect 116801 157961 116829 157989
rect 132099 158147 132127 158175
rect 132161 158147 132189 158175
rect 132099 158085 132127 158113
rect 132161 158085 132189 158113
rect 132099 158023 132127 158051
rect 132161 158023 132189 158051
rect 132099 157961 132127 157989
rect 132161 157961 132189 157989
rect 147459 158147 147487 158175
rect 147521 158147 147549 158175
rect 147459 158085 147487 158113
rect 147521 158085 147549 158113
rect 147459 158023 147487 158051
rect 147521 158023 147549 158051
rect 147459 157961 147487 157989
rect 147521 157961 147549 157989
rect 162819 158147 162847 158175
rect 162881 158147 162909 158175
rect 162819 158085 162847 158113
rect 162881 158085 162909 158113
rect 162819 158023 162847 158051
rect 162881 158023 162909 158051
rect 162819 157961 162847 157989
rect 162881 157961 162909 157989
rect 178179 158147 178207 158175
rect 178241 158147 178269 158175
rect 178179 158085 178207 158113
rect 178241 158085 178269 158113
rect 178179 158023 178207 158051
rect 178241 158023 178269 158051
rect 178179 157961 178207 157989
rect 178241 157961 178269 157989
rect 193539 158147 193567 158175
rect 193601 158147 193629 158175
rect 193539 158085 193567 158113
rect 193601 158085 193629 158113
rect 193539 158023 193567 158051
rect 193601 158023 193629 158051
rect 193539 157961 193567 157989
rect 193601 157961 193629 157989
rect 217797 298578 217825 298606
rect 217859 298578 217887 298606
rect 217921 298578 217949 298606
rect 217983 298578 218011 298606
rect 217797 298516 217825 298544
rect 217859 298516 217887 298544
rect 217921 298516 217949 298544
rect 217983 298516 218011 298544
rect 217797 298454 217825 298482
rect 217859 298454 217887 298482
rect 217921 298454 217949 298482
rect 217983 298454 218011 298482
rect 217797 298392 217825 298420
rect 217859 298392 217887 298420
rect 217921 298392 217949 298420
rect 217983 298392 218011 298420
rect 217797 290147 217825 290175
rect 217859 290147 217887 290175
rect 217921 290147 217949 290175
rect 217983 290147 218011 290175
rect 217797 290085 217825 290113
rect 217859 290085 217887 290113
rect 217921 290085 217949 290113
rect 217983 290085 218011 290113
rect 217797 290023 217825 290051
rect 217859 290023 217887 290051
rect 217921 290023 217949 290051
rect 217983 290023 218011 290051
rect 217797 289961 217825 289989
rect 217859 289961 217887 289989
rect 217921 289961 217949 289989
rect 217983 289961 218011 289989
rect 217797 281147 217825 281175
rect 217859 281147 217887 281175
rect 217921 281147 217949 281175
rect 217983 281147 218011 281175
rect 217797 281085 217825 281113
rect 217859 281085 217887 281113
rect 217921 281085 217949 281113
rect 217983 281085 218011 281113
rect 217797 281023 217825 281051
rect 217859 281023 217887 281051
rect 217921 281023 217949 281051
rect 217983 281023 218011 281051
rect 217797 280961 217825 280989
rect 217859 280961 217887 280989
rect 217921 280961 217949 280989
rect 217983 280961 218011 280989
rect 217797 272147 217825 272175
rect 217859 272147 217887 272175
rect 217921 272147 217949 272175
rect 217983 272147 218011 272175
rect 217797 272085 217825 272113
rect 217859 272085 217887 272113
rect 217921 272085 217949 272113
rect 217983 272085 218011 272113
rect 217797 272023 217825 272051
rect 217859 272023 217887 272051
rect 217921 272023 217949 272051
rect 217983 272023 218011 272051
rect 217797 271961 217825 271989
rect 217859 271961 217887 271989
rect 217921 271961 217949 271989
rect 217983 271961 218011 271989
rect 217797 263147 217825 263175
rect 217859 263147 217887 263175
rect 217921 263147 217949 263175
rect 217983 263147 218011 263175
rect 217797 263085 217825 263113
rect 217859 263085 217887 263113
rect 217921 263085 217949 263113
rect 217983 263085 218011 263113
rect 217797 263023 217825 263051
rect 217859 263023 217887 263051
rect 217921 263023 217949 263051
rect 217983 263023 218011 263051
rect 217797 262961 217825 262989
rect 217859 262961 217887 262989
rect 217921 262961 217949 262989
rect 217983 262961 218011 262989
rect 217797 254147 217825 254175
rect 217859 254147 217887 254175
rect 217921 254147 217949 254175
rect 217983 254147 218011 254175
rect 217797 254085 217825 254113
rect 217859 254085 217887 254113
rect 217921 254085 217949 254113
rect 217983 254085 218011 254113
rect 217797 254023 217825 254051
rect 217859 254023 217887 254051
rect 217921 254023 217949 254051
rect 217983 254023 218011 254051
rect 217797 253961 217825 253989
rect 217859 253961 217887 253989
rect 217921 253961 217949 253989
rect 217983 253961 218011 253989
rect 217797 245147 217825 245175
rect 217859 245147 217887 245175
rect 217921 245147 217949 245175
rect 217983 245147 218011 245175
rect 217797 245085 217825 245113
rect 217859 245085 217887 245113
rect 217921 245085 217949 245113
rect 217983 245085 218011 245113
rect 217797 245023 217825 245051
rect 217859 245023 217887 245051
rect 217921 245023 217949 245051
rect 217983 245023 218011 245051
rect 217797 244961 217825 244989
rect 217859 244961 217887 244989
rect 217921 244961 217949 244989
rect 217983 244961 218011 244989
rect 217797 236147 217825 236175
rect 217859 236147 217887 236175
rect 217921 236147 217949 236175
rect 217983 236147 218011 236175
rect 217797 236085 217825 236113
rect 217859 236085 217887 236113
rect 217921 236085 217949 236113
rect 217983 236085 218011 236113
rect 217797 236023 217825 236051
rect 217859 236023 217887 236051
rect 217921 236023 217949 236051
rect 217983 236023 218011 236051
rect 217797 235961 217825 235989
rect 217859 235961 217887 235989
rect 217921 235961 217949 235989
rect 217983 235961 218011 235989
rect 217797 227147 217825 227175
rect 217859 227147 217887 227175
rect 217921 227147 217949 227175
rect 217983 227147 218011 227175
rect 217797 227085 217825 227113
rect 217859 227085 217887 227113
rect 217921 227085 217949 227113
rect 217983 227085 218011 227113
rect 217797 227023 217825 227051
rect 217859 227023 217887 227051
rect 217921 227023 217949 227051
rect 217983 227023 218011 227051
rect 217797 226961 217825 226989
rect 217859 226961 217887 226989
rect 217921 226961 217949 226989
rect 217983 226961 218011 226989
rect 217797 218147 217825 218175
rect 217859 218147 217887 218175
rect 217921 218147 217949 218175
rect 217983 218147 218011 218175
rect 217797 218085 217825 218113
rect 217859 218085 217887 218113
rect 217921 218085 217949 218113
rect 217983 218085 218011 218113
rect 217797 218023 217825 218051
rect 217859 218023 217887 218051
rect 217921 218023 217949 218051
rect 217983 218023 218011 218051
rect 217797 217961 217825 217989
rect 217859 217961 217887 217989
rect 217921 217961 217949 217989
rect 217983 217961 218011 217989
rect 217797 209147 217825 209175
rect 217859 209147 217887 209175
rect 217921 209147 217949 209175
rect 217983 209147 218011 209175
rect 217797 209085 217825 209113
rect 217859 209085 217887 209113
rect 217921 209085 217949 209113
rect 217983 209085 218011 209113
rect 217797 209023 217825 209051
rect 217859 209023 217887 209051
rect 217921 209023 217949 209051
rect 217983 209023 218011 209051
rect 217797 208961 217825 208989
rect 217859 208961 217887 208989
rect 217921 208961 217949 208989
rect 217983 208961 218011 208989
rect 217797 200147 217825 200175
rect 217859 200147 217887 200175
rect 217921 200147 217949 200175
rect 217983 200147 218011 200175
rect 217797 200085 217825 200113
rect 217859 200085 217887 200113
rect 217921 200085 217949 200113
rect 217983 200085 218011 200113
rect 217797 200023 217825 200051
rect 217859 200023 217887 200051
rect 217921 200023 217949 200051
rect 217983 200023 218011 200051
rect 217797 199961 217825 199989
rect 217859 199961 217887 199989
rect 217921 199961 217949 199989
rect 217983 199961 218011 199989
rect 217797 191147 217825 191175
rect 217859 191147 217887 191175
rect 217921 191147 217949 191175
rect 217983 191147 218011 191175
rect 217797 191085 217825 191113
rect 217859 191085 217887 191113
rect 217921 191085 217949 191113
rect 217983 191085 218011 191113
rect 217797 191023 217825 191051
rect 217859 191023 217887 191051
rect 217921 191023 217949 191051
rect 217983 191023 218011 191051
rect 217797 190961 217825 190989
rect 217859 190961 217887 190989
rect 217921 190961 217949 190989
rect 217983 190961 218011 190989
rect 217797 182147 217825 182175
rect 217859 182147 217887 182175
rect 217921 182147 217949 182175
rect 217983 182147 218011 182175
rect 217797 182085 217825 182113
rect 217859 182085 217887 182113
rect 217921 182085 217949 182113
rect 217983 182085 218011 182113
rect 217797 182023 217825 182051
rect 217859 182023 217887 182051
rect 217921 182023 217949 182051
rect 217983 182023 218011 182051
rect 217797 181961 217825 181989
rect 217859 181961 217887 181989
rect 217921 181961 217949 181989
rect 217983 181961 218011 181989
rect 217797 173147 217825 173175
rect 217859 173147 217887 173175
rect 217921 173147 217949 173175
rect 217983 173147 218011 173175
rect 217797 173085 217825 173113
rect 217859 173085 217887 173113
rect 217921 173085 217949 173113
rect 217983 173085 218011 173113
rect 217797 173023 217825 173051
rect 217859 173023 217887 173051
rect 217921 173023 217949 173051
rect 217983 173023 218011 173051
rect 217797 172961 217825 172989
rect 217859 172961 217887 172989
rect 217921 172961 217949 172989
rect 217983 172961 218011 172989
rect 217797 164147 217825 164175
rect 217859 164147 217887 164175
rect 217921 164147 217949 164175
rect 217983 164147 218011 164175
rect 217797 164085 217825 164113
rect 217859 164085 217887 164113
rect 217921 164085 217949 164113
rect 217983 164085 218011 164113
rect 217797 164023 217825 164051
rect 217859 164023 217887 164051
rect 217921 164023 217949 164051
rect 217983 164023 218011 164051
rect 217797 163961 217825 163989
rect 217859 163961 217887 163989
rect 217921 163961 217949 163989
rect 217983 163961 218011 163989
rect 204297 158147 204325 158175
rect 204359 158147 204387 158175
rect 204421 158147 204449 158175
rect 204483 158147 204511 158175
rect 204297 158085 204325 158113
rect 204359 158085 204387 158113
rect 204421 158085 204449 158113
rect 204483 158085 204511 158113
rect 204297 158023 204325 158051
rect 204359 158023 204387 158051
rect 204421 158023 204449 158051
rect 204483 158023 204511 158051
rect 204297 157961 204325 157989
rect 204359 157961 204387 157989
rect 204421 157961 204449 157989
rect 204483 157961 204511 157989
rect 109059 155147 109087 155175
rect 109121 155147 109149 155175
rect 109059 155085 109087 155113
rect 109121 155085 109149 155113
rect 109059 155023 109087 155051
rect 109121 155023 109149 155051
rect 109059 154961 109087 154989
rect 109121 154961 109149 154989
rect 124419 155147 124447 155175
rect 124481 155147 124509 155175
rect 124419 155085 124447 155113
rect 124481 155085 124509 155113
rect 124419 155023 124447 155051
rect 124481 155023 124509 155051
rect 124419 154961 124447 154989
rect 124481 154961 124509 154989
rect 139779 155147 139807 155175
rect 139841 155147 139869 155175
rect 139779 155085 139807 155113
rect 139841 155085 139869 155113
rect 139779 155023 139807 155051
rect 139841 155023 139869 155051
rect 139779 154961 139807 154989
rect 139841 154961 139869 154989
rect 155139 155147 155167 155175
rect 155201 155147 155229 155175
rect 155139 155085 155167 155113
rect 155201 155085 155229 155113
rect 155139 155023 155167 155051
rect 155201 155023 155229 155051
rect 155139 154961 155167 154989
rect 155201 154961 155229 154989
rect 170499 155147 170527 155175
rect 170561 155147 170589 155175
rect 170499 155085 170527 155113
rect 170561 155085 170589 155113
rect 170499 155023 170527 155051
rect 170561 155023 170589 155051
rect 170499 154961 170527 154989
rect 170561 154961 170589 154989
rect 185859 155147 185887 155175
rect 185921 155147 185949 155175
rect 185859 155085 185887 155113
rect 185921 155085 185949 155113
rect 185859 155023 185887 155051
rect 185921 155023 185949 155051
rect 185859 154961 185887 154989
rect 185921 154961 185949 154989
rect 201219 155147 201247 155175
rect 201281 155147 201309 155175
rect 201219 155085 201247 155113
rect 201281 155085 201309 155113
rect 201219 155023 201247 155051
rect 201281 155023 201309 155051
rect 201219 154961 201247 154989
rect 201281 154961 201309 154989
rect 96777 149147 96805 149175
rect 96839 149147 96867 149175
rect 96901 149147 96929 149175
rect 96963 149147 96991 149175
rect 96777 149085 96805 149113
rect 96839 149085 96867 149113
rect 96901 149085 96929 149113
rect 96963 149085 96991 149113
rect 96777 149023 96805 149051
rect 96839 149023 96867 149051
rect 96901 149023 96929 149051
rect 96963 149023 96991 149051
rect 96777 148961 96805 148989
rect 96839 148961 96867 148989
rect 96901 148961 96929 148989
rect 96963 148961 96991 148989
rect 101379 149147 101407 149175
rect 101441 149147 101469 149175
rect 101379 149085 101407 149113
rect 101441 149085 101469 149113
rect 101379 149023 101407 149051
rect 101441 149023 101469 149051
rect 101379 148961 101407 148989
rect 101441 148961 101469 148989
rect 116739 149147 116767 149175
rect 116801 149147 116829 149175
rect 116739 149085 116767 149113
rect 116801 149085 116829 149113
rect 116739 149023 116767 149051
rect 116801 149023 116829 149051
rect 116739 148961 116767 148989
rect 116801 148961 116829 148989
rect 132099 149147 132127 149175
rect 132161 149147 132189 149175
rect 132099 149085 132127 149113
rect 132161 149085 132189 149113
rect 132099 149023 132127 149051
rect 132161 149023 132189 149051
rect 132099 148961 132127 148989
rect 132161 148961 132189 148989
rect 147459 149147 147487 149175
rect 147521 149147 147549 149175
rect 147459 149085 147487 149113
rect 147521 149085 147549 149113
rect 147459 149023 147487 149051
rect 147521 149023 147549 149051
rect 147459 148961 147487 148989
rect 147521 148961 147549 148989
rect 162819 149147 162847 149175
rect 162881 149147 162909 149175
rect 162819 149085 162847 149113
rect 162881 149085 162909 149113
rect 162819 149023 162847 149051
rect 162881 149023 162909 149051
rect 162819 148961 162847 148989
rect 162881 148961 162909 148989
rect 178179 149147 178207 149175
rect 178241 149147 178269 149175
rect 178179 149085 178207 149113
rect 178241 149085 178269 149113
rect 178179 149023 178207 149051
rect 178241 149023 178269 149051
rect 178179 148961 178207 148989
rect 178241 148961 178269 148989
rect 193539 149147 193567 149175
rect 193601 149147 193629 149175
rect 193539 149085 193567 149113
rect 193601 149085 193629 149113
rect 193539 149023 193567 149051
rect 193601 149023 193629 149051
rect 193539 148961 193567 148989
rect 193601 148961 193629 148989
rect 208899 158147 208927 158175
rect 208961 158147 208989 158175
rect 208899 158085 208927 158113
rect 208961 158085 208989 158113
rect 208899 158023 208927 158051
rect 208961 158023 208989 158051
rect 208899 157961 208927 157989
rect 208961 157961 208989 157989
rect 216579 155147 216607 155175
rect 216641 155147 216669 155175
rect 216579 155085 216607 155113
rect 216641 155085 216669 155113
rect 216579 155023 216607 155051
rect 216641 155023 216669 155051
rect 216579 154961 216607 154989
rect 216641 154961 216669 154989
rect 217797 155147 217825 155175
rect 217859 155147 217887 155175
rect 217921 155147 217949 155175
rect 217983 155147 218011 155175
rect 217797 155085 217825 155113
rect 217859 155085 217887 155113
rect 217921 155085 217949 155113
rect 217983 155085 218011 155113
rect 217797 155023 217825 155051
rect 217859 155023 217887 155051
rect 217921 155023 217949 155051
rect 217983 155023 218011 155051
rect 217797 154961 217825 154989
rect 217859 154961 217887 154989
rect 217921 154961 217949 154989
rect 217983 154961 218011 154989
rect 204297 149147 204325 149175
rect 204359 149147 204387 149175
rect 204421 149147 204449 149175
rect 204483 149147 204511 149175
rect 204297 149085 204325 149113
rect 204359 149085 204387 149113
rect 204421 149085 204449 149113
rect 204483 149085 204511 149113
rect 204297 149023 204325 149051
rect 204359 149023 204387 149051
rect 204421 149023 204449 149051
rect 204483 149023 204511 149051
rect 204297 148961 204325 148989
rect 204359 148961 204387 148989
rect 204421 148961 204449 148989
rect 204483 148961 204511 148989
rect 109059 146147 109087 146175
rect 109121 146147 109149 146175
rect 109059 146085 109087 146113
rect 109121 146085 109149 146113
rect 109059 146023 109087 146051
rect 109121 146023 109149 146051
rect 109059 145961 109087 145989
rect 109121 145961 109149 145989
rect 124419 146147 124447 146175
rect 124481 146147 124509 146175
rect 124419 146085 124447 146113
rect 124481 146085 124509 146113
rect 124419 146023 124447 146051
rect 124481 146023 124509 146051
rect 124419 145961 124447 145989
rect 124481 145961 124509 145989
rect 139779 146147 139807 146175
rect 139841 146147 139869 146175
rect 139779 146085 139807 146113
rect 139841 146085 139869 146113
rect 139779 146023 139807 146051
rect 139841 146023 139869 146051
rect 139779 145961 139807 145989
rect 139841 145961 139869 145989
rect 155139 146147 155167 146175
rect 155201 146147 155229 146175
rect 155139 146085 155167 146113
rect 155201 146085 155229 146113
rect 155139 146023 155167 146051
rect 155201 146023 155229 146051
rect 155139 145961 155167 145989
rect 155201 145961 155229 145989
rect 170499 146147 170527 146175
rect 170561 146147 170589 146175
rect 170499 146085 170527 146113
rect 170561 146085 170589 146113
rect 170499 146023 170527 146051
rect 170561 146023 170589 146051
rect 170499 145961 170527 145989
rect 170561 145961 170589 145989
rect 185859 146147 185887 146175
rect 185921 146147 185949 146175
rect 185859 146085 185887 146113
rect 185921 146085 185949 146113
rect 185859 146023 185887 146051
rect 185921 146023 185949 146051
rect 185859 145961 185887 145989
rect 185921 145961 185949 145989
rect 201219 146147 201247 146175
rect 201281 146147 201309 146175
rect 201219 146085 201247 146113
rect 201281 146085 201309 146113
rect 201219 146023 201247 146051
rect 201281 146023 201309 146051
rect 201219 145961 201247 145989
rect 201281 145961 201309 145989
rect 96777 140147 96805 140175
rect 96839 140147 96867 140175
rect 96901 140147 96929 140175
rect 96963 140147 96991 140175
rect 96777 140085 96805 140113
rect 96839 140085 96867 140113
rect 96901 140085 96929 140113
rect 96963 140085 96991 140113
rect 96777 140023 96805 140051
rect 96839 140023 96867 140051
rect 96901 140023 96929 140051
rect 96963 140023 96991 140051
rect 96777 139961 96805 139989
rect 96839 139961 96867 139989
rect 96901 139961 96929 139989
rect 96963 139961 96991 139989
rect 101379 140147 101407 140175
rect 101441 140147 101469 140175
rect 101379 140085 101407 140113
rect 101441 140085 101469 140113
rect 101379 140023 101407 140051
rect 101441 140023 101469 140051
rect 101379 139961 101407 139989
rect 101441 139961 101469 139989
rect 116739 140147 116767 140175
rect 116801 140147 116829 140175
rect 116739 140085 116767 140113
rect 116801 140085 116829 140113
rect 116739 140023 116767 140051
rect 116801 140023 116829 140051
rect 116739 139961 116767 139989
rect 116801 139961 116829 139989
rect 132099 140147 132127 140175
rect 132161 140147 132189 140175
rect 132099 140085 132127 140113
rect 132161 140085 132189 140113
rect 132099 140023 132127 140051
rect 132161 140023 132189 140051
rect 132099 139961 132127 139989
rect 132161 139961 132189 139989
rect 147459 140147 147487 140175
rect 147521 140147 147549 140175
rect 147459 140085 147487 140113
rect 147521 140085 147549 140113
rect 147459 140023 147487 140051
rect 147521 140023 147549 140051
rect 147459 139961 147487 139989
rect 147521 139961 147549 139989
rect 162819 140147 162847 140175
rect 162881 140147 162909 140175
rect 162819 140085 162847 140113
rect 162881 140085 162909 140113
rect 162819 140023 162847 140051
rect 162881 140023 162909 140051
rect 162819 139961 162847 139989
rect 162881 139961 162909 139989
rect 178179 140147 178207 140175
rect 178241 140147 178269 140175
rect 178179 140085 178207 140113
rect 178241 140085 178269 140113
rect 178179 140023 178207 140051
rect 178241 140023 178269 140051
rect 178179 139961 178207 139989
rect 178241 139961 178269 139989
rect 193539 140147 193567 140175
rect 193601 140147 193629 140175
rect 193539 140085 193567 140113
rect 193601 140085 193629 140113
rect 193539 140023 193567 140051
rect 193601 140023 193629 140051
rect 193539 139961 193567 139989
rect 193601 139961 193629 139989
rect 208899 149147 208927 149175
rect 208961 149147 208989 149175
rect 208899 149085 208927 149113
rect 208961 149085 208989 149113
rect 208899 149023 208927 149051
rect 208961 149023 208989 149051
rect 208899 148961 208927 148989
rect 208961 148961 208989 148989
rect 216579 146147 216607 146175
rect 216641 146147 216669 146175
rect 216579 146085 216607 146113
rect 216641 146085 216669 146113
rect 216579 146023 216607 146051
rect 216641 146023 216669 146051
rect 216579 145961 216607 145989
rect 216641 145961 216669 145989
rect 217797 146147 217825 146175
rect 217859 146147 217887 146175
rect 217921 146147 217949 146175
rect 217983 146147 218011 146175
rect 217797 146085 217825 146113
rect 217859 146085 217887 146113
rect 217921 146085 217949 146113
rect 217983 146085 218011 146113
rect 217797 146023 217825 146051
rect 217859 146023 217887 146051
rect 217921 146023 217949 146051
rect 217983 146023 218011 146051
rect 217797 145961 217825 145989
rect 217859 145961 217887 145989
rect 217921 145961 217949 145989
rect 217983 145961 218011 145989
rect 204297 140147 204325 140175
rect 204359 140147 204387 140175
rect 204421 140147 204449 140175
rect 204483 140147 204511 140175
rect 204297 140085 204325 140113
rect 204359 140085 204387 140113
rect 204421 140085 204449 140113
rect 204483 140085 204511 140113
rect 204297 140023 204325 140051
rect 204359 140023 204387 140051
rect 204421 140023 204449 140051
rect 204483 140023 204511 140051
rect 204297 139961 204325 139989
rect 204359 139961 204387 139989
rect 204421 139961 204449 139989
rect 204483 139961 204511 139989
rect 109059 137147 109087 137175
rect 109121 137147 109149 137175
rect 109059 137085 109087 137113
rect 109121 137085 109149 137113
rect 109059 137023 109087 137051
rect 109121 137023 109149 137051
rect 109059 136961 109087 136989
rect 109121 136961 109149 136989
rect 124419 137147 124447 137175
rect 124481 137147 124509 137175
rect 124419 137085 124447 137113
rect 124481 137085 124509 137113
rect 124419 137023 124447 137051
rect 124481 137023 124509 137051
rect 124419 136961 124447 136989
rect 124481 136961 124509 136989
rect 139779 137147 139807 137175
rect 139841 137147 139869 137175
rect 139779 137085 139807 137113
rect 139841 137085 139869 137113
rect 139779 137023 139807 137051
rect 139841 137023 139869 137051
rect 139779 136961 139807 136989
rect 139841 136961 139869 136989
rect 155139 137147 155167 137175
rect 155201 137147 155229 137175
rect 155139 137085 155167 137113
rect 155201 137085 155229 137113
rect 155139 137023 155167 137051
rect 155201 137023 155229 137051
rect 155139 136961 155167 136989
rect 155201 136961 155229 136989
rect 170499 137147 170527 137175
rect 170561 137147 170589 137175
rect 170499 137085 170527 137113
rect 170561 137085 170589 137113
rect 170499 137023 170527 137051
rect 170561 137023 170589 137051
rect 170499 136961 170527 136989
rect 170561 136961 170589 136989
rect 185859 137147 185887 137175
rect 185921 137147 185949 137175
rect 185859 137085 185887 137113
rect 185921 137085 185949 137113
rect 185859 137023 185887 137051
rect 185921 137023 185949 137051
rect 185859 136961 185887 136989
rect 185921 136961 185949 136989
rect 201219 137147 201247 137175
rect 201281 137147 201309 137175
rect 201219 137085 201247 137113
rect 201281 137085 201309 137113
rect 201219 137023 201247 137051
rect 201281 137023 201309 137051
rect 201219 136961 201247 136989
rect 201281 136961 201309 136989
rect 96777 131147 96805 131175
rect 96839 131147 96867 131175
rect 96901 131147 96929 131175
rect 96963 131147 96991 131175
rect 96777 131085 96805 131113
rect 96839 131085 96867 131113
rect 96901 131085 96929 131113
rect 96963 131085 96991 131113
rect 96777 131023 96805 131051
rect 96839 131023 96867 131051
rect 96901 131023 96929 131051
rect 96963 131023 96991 131051
rect 208899 140147 208927 140175
rect 208961 140147 208989 140175
rect 208899 140085 208927 140113
rect 208961 140085 208989 140113
rect 208899 140023 208927 140051
rect 208961 140023 208989 140051
rect 208899 139961 208927 139989
rect 208961 139961 208989 139989
rect 216579 137147 216607 137175
rect 216641 137147 216669 137175
rect 216579 137085 216607 137113
rect 216641 137085 216669 137113
rect 216579 137023 216607 137051
rect 216641 137023 216669 137051
rect 216579 136961 216607 136989
rect 216641 136961 216669 136989
rect 217797 137147 217825 137175
rect 217859 137147 217887 137175
rect 217921 137147 217949 137175
rect 217983 137147 218011 137175
rect 217797 137085 217825 137113
rect 217859 137085 217887 137113
rect 217921 137085 217949 137113
rect 217983 137085 218011 137113
rect 217797 137023 217825 137051
rect 217859 137023 217887 137051
rect 217921 137023 217949 137051
rect 217983 137023 218011 137051
rect 217797 136961 217825 136989
rect 217859 136961 217887 136989
rect 217921 136961 217949 136989
rect 217983 136961 218011 136989
rect 204297 131147 204325 131175
rect 204359 131147 204387 131175
rect 204421 131147 204449 131175
rect 204483 131147 204511 131175
rect 204297 131085 204325 131113
rect 204359 131085 204387 131113
rect 204421 131085 204449 131113
rect 204483 131085 204511 131113
rect 96777 130961 96805 130989
rect 96839 130961 96867 130989
rect 96901 130961 96929 130989
rect 96963 130961 96991 130989
rect 112137 130986 112165 131014
rect 112199 130986 112227 131014
rect 112261 130986 112289 131014
rect 112323 130986 112351 131014
rect 112137 130924 112165 130952
rect 112199 130924 112227 130952
rect 112261 130924 112289 130952
rect 112323 130924 112351 130952
rect 96777 122147 96805 122175
rect 96839 122147 96867 122175
rect 96901 122147 96929 122175
rect 96963 122147 96991 122175
rect 96777 122085 96805 122113
rect 96839 122085 96867 122113
rect 96901 122085 96929 122113
rect 96963 122085 96991 122113
rect 96777 122023 96805 122051
rect 96839 122023 96867 122051
rect 96901 122023 96929 122051
rect 96963 122023 96991 122051
rect 96777 121961 96805 121989
rect 96839 121961 96867 121989
rect 96901 121961 96929 121989
rect 96963 121961 96991 121989
rect 109939 122147 109967 122175
rect 110001 122147 110029 122175
rect 109939 122085 109967 122113
rect 110001 122085 110029 122113
rect 109939 122023 109967 122051
rect 110001 122023 110029 122051
rect 109939 121961 109967 121989
rect 110001 121961 110029 121989
rect 125637 128147 125665 128175
rect 125699 128147 125727 128175
rect 125761 128147 125789 128175
rect 125823 128147 125851 128175
rect 125637 128085 125665 128113
rect 125699 128085 125727 128113
rect 125761 128085 125789 128113
rect 125823 128085 125851 128113
rect 125637 128023 125665 128051
rect 125699 128023 125727 128051
rect 125761 128023 125789 128051
rect 125823 128023 125851 128051
rect 125637 127961 125665 127989
rect 125699 127961 125727 127989
rect 125761 127961 125789 127989
rect 125823 127961 125851 127989
rect 112137 122147 112165 122175
rect 112199 122147 112227 122175
rect 112261 122147 112289 122175
rect 112323 122147 112351 122175
rect 112137 122085 112165 122113
rect 112199 122085 112227 122113
rect 112261 122085 112289 122113
rect 112323 122085 112351 122113
rect 112137 122023 112165 122051
rect 112199 122023 112227 122051
rect 112261 122023 112289 122051
rect 112323 122023 112351 122051
rect 112137 121961 112165 121989
rect 112199 121961 112227 121989
rect 112261 121961 112289 121989
rect 112323 121961 112351 121989
rect 125299 122147 125327 122175
rect 125361 122147 125389 122175
rect 125299 122085 125327 122113
rect 125361 122085 125389 122113
rect 125299 122023 125327 122051
rect 125361 122023 125389 122051
rect 125299 121961 125327 121989
rect 125361 121961 125389 121989
rect 102259 119147 102287 119175
rect 102321 119147 102349 119175
rect 102259 119085 102287 119113
rect 102321 119085 102349 119113
rect 102259 119023 102287 119051
rect 102321 119023 102349 119051
rect 102259 118961 102287 118989
rect 102321 118961 102349 118989
rect 117619 119147 117647 119175
rect 117681 119147 117709 119175
rect 117619 119085 117647 119113
rect 117681 119085 117709 119113
rect 117619 119023 117647 119051
rect 117681 119023 117709 119051
rect 117619 118961 117647 118989
rect 117681 118961 117709 118989
rect 125637 119147 125665 119175
rect 125699 119147 125727 119175
rect 125761 119147 125789 119175
rect 125823 119147 125851 119175
rect 125637 119085 125665 119113
rect 125699 119085 125727 119113
rect 125761 119085 125789 119113
rect 125823 119085 125851 119113
rect 125637 119023 125665 119051
rect 125699 119023 125727 119051
rect 125761 119023 125789 119051
rect 125823 119023 125851 119051
rect 125637 118961 125665 118989
rect 125699 118961 125727 118989
rect 125761 118961 125789 118989
rect 125823 118961 125851 118989
rect 96777 113147 96805 113175
rect 96839 113147 96867 113175
rect 96901 113147 96929 113175
rect 96963 113147 96991 113175
rect 96777 113085 96805 113113
rect 96839 113085 96867 113113
rect 96901 113085 96929 113113
rect 96963 113085 96991 113113
rect 96777 113023 96805 113051
rect 96839 113023 96867 113051
rect 96901 113023 96929 113051
rect 96963 113023 96991 113051
rect 96777 112961 96805 112989
rect 96839 112961 96867 112989
rect 96901 112961 96929 112989
rect 96963 112961 96991 112989
rect 109939 113147 109967 113175
rect 110001 113147 110029 113175
rect 109939 113085 109967 113113
rect 110001 113085 110029 113113
rect 109939 113023 109967 113051
rect 110001 113023 110029 113051
rect 109939 112961 109967 112989
rect 110001 112961 110029 112989
rect 125299 113147 125327 113175
rect 125361 113147 125389 113175
rect 125299 113085 125327 113113
rect 125361 113085 125389 113113
rect 125299 113023 125327 113051
rect 125361 113023 125389 113051
rect 125299 112961 125327 112989
rect 125361 112961 125389 112989
rect 102259 110147 102287 110175
rect 102321 110147 102349 110175
rect 102259 110085 102287 110113
rect 102321 110085 102349 110113
rect 102259 110023 102287 110051
rect 102321 110023 102349 110051
rect 102259 109961 102287 109989
rect 102321 109961 102349 109989
rect 117619 110147 117647 110175
rect 117681 110147 117709 110175
rect 117619 110085 117647 110113
rect 117681 110085 117709 110113
rect 117619 110023 117647 110051
rect 117681 110023 117709 110051
rect 117619 109961 117647 109989
rect 117681 109961 117709 109989
rect 125637 110147 125665 110175
rect 125699 110147 125727 110175
rect 125761 110147 125789 110175
rect 125823 110147 125851 110175
rect 125637 110085 125665 110113
rect 125699 110085 125727 110113
rect 125761 110085 125789 110113
rect 125823 110085 125851 110113
rect 125637 110023 125665 110051
rect 125699 110023 125727 110051
rect 125761 110023 125789 110051
rect 125823 110023 125851 110051
rect 125637 109961 125665 109989
rect 125699 109961 125727 109989
rect 125761 109961 125789 109989
rect 125823 109961 125851 109989
rect 96777 104147 96805 104175
rect 96839 104147 96867 104175
rect 96901 104147 96929 104175
rect 96963 104147 96991 104175
rect 96777 104085 96805 104113
rect 96839 104085 96867 104113
rect 96901 104085 96929 104113
rect 96963 104085 96991 104113
rect 96777 104023 96805 104051
rect 96839 104023 96867 104051
rect 96901 104023 96929 104051
rect 96963 104023 96991 104051
rect 96777 103961 96805 103989
rect 96839 103961 96867 103989
rect 96901 103961 96929 103989
rect 96963 103961 96991 103989
rect 109939 104147 109967 104175
rect 110001 104147 110029 104175
rect 109939 104085 109967 104113
rect 110001 104085 110029 104113
rect 109939 104023 109967 104051
rect 110001 104023 110029 104051
rect 109939 103961 109967 103989
rect 110001 103961 110029 103989
rect 125299 104147 125327 104175
rect 125361 104147 125389 104175
rect 125299 104085 125327 104113
rect 125361 104085 125389 104113
rect 125299 104023 125327 104051
rect 125361 104023 125389 104051
rect 125299 103961 125327 103989
rect 125361 103961 125389 103989
rect 102259 101147 102287 101175
rect 102321 101147 102349 101175
rect 102259 101085 102287 101113
rect 102321 101085 102349 101113
rect 102259 101023 102287 101051
rect 102321 101023 102349 101051
rect 102259 100961 102287 100989
rect 102321 100961 102349 100989
rect 117619 101147 117647 101175
rect 117681 101147 117709 101175
rect 117619 101085 117647 101113
rect 117681 101085 117709 101113
rect 117619 101023 117647 101051
rect 117681 101023 117709 101051
rect 117619 100961 117647 100989
rect 117681 100961 117709 100989
rect 125637 101147 125665 101175
rect 125699 101147 125727 101175
rect 125761 101147 125789 101175
rect 125823 101147 125851 101175
rect 125637 101085 125665 101113
rect 125699 101085 125727 101113
rect 125761 101085 125789 101113
rect 125823 101085 125851 101113
rect 125637 101023 125665 101051
rect 125699 101023 125727 101051
rect 125761 101023 125789 101051
rect 125823 101023 125851 101051
rect 125637 100961 125665 100989
rect 125699 100961 125727 100989
rect 125761 100961 125789 100989
rect 125823 100961 125851 100989
rect 96777 95147 96805 95175
rect 96839 95147 96867 95175
rect 96901 95147 96929 95175
rect 96963 95147 96991 95175
rect 96777 95085 96805 95113
rect 96839 95085 96867 95113
rect 96901 95085 96929 95113
rect 96963 95085 96991 95113
rect 96777 95023 96805 95051
rect 96839 95023 96867 95051
rect 96901 95023 96929 95051
rect 96963 95023 96991 95051
rect 96777 94961 96805 94989
rect 96839 94961 96867 94989
rect 96901 94961 96929 94989
rect 96963 94961 96991 94989
rect 96777 86147 96805 86175
rect 96839 86147 96867 86175
rect 96901 86147 96929 86175
rect 96963 86147 96991 86175
rect 96777 86085 96805 86113
rect 96839 86085 96867 86113
rect 96901 86085 96929 86113
rect 96963 86085 96991 86113
rect 96777 86023 96805 86051
rect 96839 86023 96867 86051
rect 96901 86023 96929 86051
rect 96963 86023 96991 86051
rect 96777 85961 96805 85989
rect 96839 85961 96867 85989
rect 96901 85961 96929 85989
rect 96963 85961 96991 85989
rect 96777 77147 96805 77175
rect 96839 77147 96867 77175
rect 96901 77147 96929 77175
rect 96963 77147 96991 77175
rect 96777 77085 96805 77113
rect 96839 77085 96867 77113
rect 96901 77085 96929 77113
rect 96963 77085 96991 77113
rect 96777 77023 96805 77051
rect 96839 77023 96867 77051
rect 96901 77023 96929 77051
rect 96963 77023 96991 77051
rect 96777 76961 96805 76989
rect 96839 76961 96867 76989
rect 96901 76961 96929 76989
rect 96963 76961 96991 76989
rect 96777 68147 96805 68175
rect 96839 68147 96867 68175
rect 96901 68147 96929 68175
rect 96963 68147 96991 68175
rect 96777 68085 96805 68113
rect 96839 68085 96867 68113
rect 96901 68085 96929 68113
rect 96963 68085 96991 68113
rect 96777 68023 96805 68051
rect 96839 68023 96867 68051
rect 96901 68023 96929 68051
rect 96963 68023 96991 68051
rect 96777 67961 96805 67989
rect 96839 67961 96867 67989
rect 96901 67961 96929 67989
rect 96963 67961 96991 67989
rect 96777 59147 96805 59175
rect 96839 59147 96867 59175
rect 96901 59147 96929 59175
rect 96963 59147 96991 59175
rect 96777 59085 96805 59113
rect 96839 59085 96867 59113
rect 96901 59085 96929 59113
rect 96963 59085 96991 59113
rect 96777 59023 96805 59051
rect 96839 59023 96867 59051
rect 96901 59023 96929 59051
rect 96963 59023 96991 59051
rect 96777 58961 96805 58989
rect 96839 58961 96867 58989
rect 96901 58961 96929 58989
rect 96963 58961 96991 58989
rect 96777 50147 96805 50175
rect 96839 50147 96867 50175
rect 96901 50147 96929 50175
rect 96963 50147 96991 50175
rect 96777 50085 96805 50113
rect 96839 50085 96867 50113
rect 96901 50085 96929 50113
rect 96963 50085 96991 50113
rect 96777 50023 96805 50051
rect 96839 50023 96867 50051
rect 96901 50023 96929 50051
rect 96963 50023 96991 50051
rect 96777 49961 96805 49989
rect 96839 49961 96867 49989
rect 96901 49961 96929 49989
rect 96963 49961 96991 49989
rect 96777 41147 96805 41175
rect 96839 41147 96867 41175
rect 96901 41147 96929 41175
rect 96963 41147 96991 41175
rect 96777 41085 96805 41113
rect 96839 41085 96867 41113
rect 96901 41085 96929 41113
rect 96963 41085 96991 41113
rect 96777 41023 96805 41051
rect 96839 41023 96867 41051
rect 96901 41023 96929 41051
rect 96963 41023 96991 41051
rect 96777 40961 96805 40989
rect 96839 40961 96867 40989
rect 96901 40961 96929 40989
rect 96963 40961 96991 40989
rect 96777 32147 96805 32175
rect 96839 32147 96867 32175
rect 96901 32147 96929 32175
rect 96963 32147 96991 32175
rect 96777 32085 96805 32113
rect 96839 32085 96867 32113
rect 96901 32085 96929 32113
rect 96963 32085 96991 32113
rect 96777 32023 96805 32051
rect 96839 32023 96867 32051
rect 96901 32023 96929 32051
rect 96963 32023 96991 32051
rect 96777 31961 96805 31989
rect 96839 31961 96867 31989
rect 96901 31961 96929 31989
rect 96963 31961 96991 31989
rect 96777 23147 96805 23175
rect 96839 23147 96867 23175
rect 96901 23147 96929 23175
rect 96963 23147 96991 23175
rect 96777 23085 96805 23113
rect 96839 23085 96867 23113
rect 96901 23085 96929 23113
rect 96963 23085 96991 23113
rect 96777 23023 96805 23051
rect 96839 23023 96867 23051
rect 96901 23023 96929 23051
rect 96963 23023 96991 23051
rect 96777 22961 96805 22989
rect 96839 22961 96867 22989
rect 96901 22961 96929 22989
rect 96963 22961 96991 22989
rect 96777 14147 96805 14175
rect 96839 14147 96867 14175
rect 96901 14147 96929 14175
rect 96963 14147 96991 14175
rect 96777 14085 96805 14113
rect 96839 14085 96867 14113
rect 96901 14085 96929 14113
rect 96963 14085 96991 14113
rect 96777 14023 96805 14051
rect 96839 14023 96867 14051
rect 96901 14023 96929 14051
rect 96963 14023 96991 14051
rect 96777 13961 96805 13989
rect 96839 13961 96867 13989
rect 96901 13961 96929 13989
rect 96963 13961 96991 13989
rect 96777 5147 96805 5175
rect 96839 5147 96867 5175
rect 96901 5147 96929 5175
rect 96963 5147 96991 5175
rect 96777 5085 96805 5113
rect 96839 5085 96867 5113
rect 96901 5085 96929 5113
rect 96963 5085 96991 5113
rect 96777 5023 96805 5051
rect 96839 5023 96867 5051
rect 96901 5023 96929 5051
rect 96963 5023 96991 5051
rect 96777 4961 96805 4989
rect 96839 4961 96867 4989
rect 96901 4961 96929 4989
rect 96963 4961 96991 4989
rect 96777 -588 96805 -560
rect 96839 -588 96867 -560
rect 96901 -588 96929 -560
rect 96963 -588 96991 -560
rect 96777 -650 96805 -622
rect 96839 -650 96867 -622
rect 96901 -650 96929 -622
rect 96963 -650 96991 -622
rect 96777 -712 96805 -684
rect 96839 -712 96867 -684
rect 96901 -712 96929 -684
rect 96963 -712 96991 -684
rect 96777 -774 96805 -746
rect 96839 -774 96867 -746
rect 96901 -774 96929 -746
rect 96963 -774 96991 -746
rect 110277 92147 110305 92175
rect 110339 92147 110367 92175
rect 110401 92147 110429 92175
rect 110463 92147 110491 92175
rect 110277 92085 110305 92113
rect 110339 92085 110367 92113
rect 110401 92085 110429 92113
rect 110463 92085 110491 92113
rect 110277 92023 110305 92051
rect 110339 92023 110367 92051
rect 110401 92023 110429 92051
rect 110463 92023 110491 92051
rect 110277 91961 110305 91989
rect 110339 91961 110367 91989
rect 110401 91961 110429 91989
rect 110463 91961 110491 91989
rect 110277 83147 110305 83175
rect 110339 83147 110367 83175
rect 110401 83147 110429 83175
rect 110463 83147 110491 83175
rect 110277 83085 110305 83113
rect 110339 83085 110367 83113
rect 110401 83085 110429 83113
rect 110463 83085 110491 83113
rect 110277 83023 110305 83051
rect 110339 83023 110367 83051
rect 110401 83023 110429 83051
rect 110463 83023 110491 83051
rect 110277 82961 110305 82989
rect 110339 82961 110367 82989
rect 110401 82961 110429 82989
rect 110463 82961 110491 82989
rect 110277 74147 110305 74175
rect 110339 74147 110367 74175
rect 110401 74147 110429 74175
rect 110463 74147 110491 74175
rect 110277 74085 110305 74113
rect 110339 74085 110367 74113
rect 110401 74085 110429 74113
rect 110463 74085 110491 74113
rect 110277 74023 110305 74051
rect 110339 74023 110367 74051
rect 110401 74023 110429 74051
rect 110463 74023 110491 74051
rect 110277 73961 110305 73989
rect 110339 73961 110367 73989
rect 110401 73961 110429 73989
rect 110463 73961 110491 73989
rect 110277 65147 110305 65175
rect 110339 65147 110367 65175
rect 110401 65147 110429 65175
rect 110463 65147 110491 65175
rect 110277 65085 110305 65113
rect 110339 65085 110367 65113
rect 110401 65085 110429 65113
rect 110463 65085 110491 65113
rect 110277 65023 110305 65051
rect 110339 65023 110367 65051
rect 110401 65023 110429 65051
rect 110463 65023 110491 65051
rect 110277 64961 110305 64989
rect 110339 64961 110367 64989
rect 110401 64961 110429 64989
rect 110463 64961 110491 64989
rect 110277 56147 110305 56175
rect 110339 56147 110367 56175
rect 110401 56147 110429 56175
rect 110463 56147 110491 56175
rect 110277 56085 110305 56113
rect 110339 56085 110367 56113
rect 110401 56085 110429 56113
rect 110463 56085 110491 56113
rect 110277 56023 110305 56051
rect 110339 56023 110367 56051
rect 110401 56023 110429 56051
rect 110463 56023 110491 56051
rect 110277 55961 110305 55989
rect 110339 55961 110367 55989
rect 110401 55961 110429 55989
rect 110463 55961 110491 55989
rect 110277 47147 110305 47175
rect 110339 47147 110367 47175
rect 110401 47147 110429 47175
rect 110463 47147 110491 47175
rect 110277 47085 110305 47113
rect 110339 47085 110367 47113
rect 110401 47085 110429 47113
rect 110463 47085 110491 47113
rect 110277 47023 110305 47051
rect 110339 47023 110367 47051
rect 110401 47023 110429 47051
rect 110463 47023 110491 47051
rect 110277 46961 110305 46989
rect 110339 46961 110367 46989
rect 110401 46961 110429 46989
rect 110463 46961 110491 46989
rect 110277 38147 110305 38175
rect 110339 38147 110367 38175
rect 110401 38147 110429 38175
rect 110463 38147 110491 38175
rect 110277 38085 110305 38113
rect 110339 38085 110367 38113
rect 110401 38085 110429 38113
rect 110463 38085 110491 38113
rect 110277 38023 110305 38051
rect 110339 38023 110367 38051
rect 110401 38023 110429 38051
rect 110463 38023 110491 38051
rect 110277 37961 110305 37989
rect 110339 37961 110367 37989
rect 110401 37961 110429 37989
rect 110463 37961 110491 37989
rect 110277 29147 110305 29175
rect 110339 29147 110367 29175
rect 110401 29147 110429 29175
rect 110463 29147 110491 29175
rect 110277 29085 110305 29113
rect 110339 29085 110367 29113
rect 110401 29085 110429 29113
rect 110463 29085 110491 29113
rect 110277 29023 110305 29051
rect 110339 29023 110367 29051
rect 110401 29023 110429 29051
rect 110463 29023 110491 29051
rect 110277 28961 110305 28989
rect 110339 28961 110367 28989
rect 110401 28961 110429 28989
rect 110463 28961 110491 28989
rect 110277 20147 110305 20175
rect 110339 20147 110367 20175
rect 110401 20147 110429 20175
rect 110463 20147 110491 20175
rect 110277 20085 110305 20113
rect 110339 20085 110367 20113
rect 110401 20085 110429 20113
rect 110463 20085 110491 20113
rect 110277 20023 110305 20051
rect 110339 20023 110367 20051
rect 110401 20023 110429 20051
rect 110463 20023 110491 20051
rect 110277 19961 110305 19989
rect 110339 19961 110367 19989
rect 110401 19961 110429 19989
rect 110463 19961 110491 19989
rect 110277 11147 110305 11175
rect 110339 11147 110367 11175
rect 110401 11147 110429 11175
rect 110463 11147 110491 11175
rect 110277 11085 110305 11113
rect 110339 11085 110367 11113
rect 110401 11085 110429 11113
rect 110463 11085 110491 11113
rect 110277 11023 110305 11051
rect 110339 11023 110367 11051
rect 110401 11023 110429 11051
rect 110463 11023 110491 11051
rect 110277 10961 110305 10989
rect 110339 10961 110367 10989
rect 110401 10961 110429 10989
rect 110463 10961 110491 10989
rect 110277 2147 110305 2175
rect 110339 2147 110367 2175
rect 110401 2147 110429 2175
rect 110463 2147 110491 2175
rect 110277 2085 110305 2113
rect 110339 2085 110367 2113
rect 110401 2085 110429 2113
rect 110463 2085 110491 2113
rect 110277 2023 110305 2051
rect 110339 2023 110367 2051
rect 110401 2023 110429 2051
rect 110463 2023 110491 2051
rect 110277 1961 110305 1989
rect 110339 1961 110367 1989
rect 110401 1961 110429 1989
rect 110463 1961 110491 1989
rect 110277 -108 110305 -80
rect 110339 -108 110367 -80
rect 110401 -108 110429 -80
rect 110463 -108 110491 -80
rect 110277 -170 110305 -142
rect 110339 -170 110367 -142
rect 110401 -170 110429 -142
rect 110463 -170 110491 -142
rect 110277 -232 110305 -204
rect 110339 -232 110367 -204
rect 110401 -232 110429 -204
rect 110463 -232 110491 -204
rect 110277 -294 110305 -266
rect 110339 -294 110367 -266
rect 110401 -294 110429 -266
rect 110463 -294 110491 -266
rect 112137 95147 112165 95175
rect 112199 95147 112227 95175
rect 112261 95147 112289 95175
rect 112323 95147 112351 95175
rect 112137 95085 112165 95113
rect 112199 95085 112227 95113
rect 112261 95085 112289 95113
rect 112323 95085 112351 95113
rect 112137 95023 112165 95051
rect 112199 95023 112227 95051
rect 112261 95023 112289 95051
rect 112323 95023 112351 95051
rect 112137 94961 112165 94989
rect 112199 94961 112227 94989
rect 112261 94961 112289 94989
rect 112323 94961 112351 94989
rect 112137 86147 112165 86175
rect 112199 86147 112227 86175
rect 112261 86147 112289 86175
rect 112323 86147 112351 86175
rect 112137 86085 112165 86113
rect 112199 86085 112227 86113
rect 112261 86085 112289 86113
rect 112323 86085 112351 86113
rect 112137 86023 112165 86051
rect 112199 86023 112227 86051
rect 112261 86023 112289 86051
rect 112323 86023 112351 86051
rect 112137 85961 112165 85989
rect 112199 85961 112227 85989
rect 112261 85961 112289 85989
rect 112323 85961 112351 85989
rect 112137 77147 112165 77175
rect 112199 77147 112227 77175
rect 112261 77147 112289 77175
rect 112323 77147 112351 77175
rect 112137 77085 112165 77113
rect 112199 77085 112227 77113
rect 112261 77085 112289 77113
rect 112323 77085 112351 77113
rect 112137 77023 112165 77051
rect 112199 77023 112227 77051
rect 112261 77023 112289 77051
rect 112323 77023 112351 77051
rect 112137 76961 112165 76989
rect 112199 76961 112227 76989
rect 112261 76961 112289 76989
rect 112323 76961 112351 76989
rect 112137 68147 112165 68175
rect 112199 68147 112227 68175
rect 112261 68147 112289 68175
rect 112323 68147 112351 68175
rect 112137 68085 112165 68113
rect 112199 68085 112227 68113
rect 112261 68085 112289 68113
rect 112323 68085 112351 68113
rect 112137 68023 112165 68051
rect 112199 68023 112227 68051
rect 112261 68023 112289 68051
rect 112323 68023 112351 68051
rect 112137 67961 112165 67989
rect 112199 67961 112227 67989
rect 112261 67961 112289 67989
rect 112323 67961 112351 67989
rect 112137 59147 112165 59175
rect 112199 59147 112227 59175
rect 112261 59147 112289 59175
rect 112323 59147 112351 59175
rect 112137 59085 112165 59113
rect 112199 59085 112227 59113
rect 112261 59085 112289 59113
rect 112323 59085 112351 59113
rect 112137 59023 112165 59051
rect 112199 59023 112227 59051
rect 112261 59023 112289 59051
rect 112323 59023 112351 59051
rect 112137 58961 112165 58989
rect 112199 58961 112227 58989
rect 112261 58961 112289 58989
rect 112323 58961 112351 58989
rect 112137 50147 112165 50175
rect 112199 50147 112227 50175
rect 112261 50147 112289 50175
rect 112323 50147 112351 50175
rect 112137 50085 112165 50113
rect 112199 50085 112227 50113
rect 112261 50085 112289 50113
rect 112323 50085 112351 50113
rect 112137 50023 112165 50051
rect 112199 50023 112227 50051
rect 112261 50023 112289 50051
rect 112323 50023 112351 50051
rect 112137 49961 112165 49989
rect 112199 49961 112227 49989
rect 112261 49961 112289 49989
rect 112323 49961 112351 49989
rect 112137 41147 112165 41175
rect 112199 41147 112227 41175
rect 112261 41147 112289 41175
rect 112323 41147 112351 41175
rect 112137 41085 112165 41113
rect 112199 41085 112227 41113
rect 112261 41085 112289 41113
rect 112323 41085 112351 41113
rect 112137 41023 112165 41051
rect 112199 41023 112227 41051
rect 112261 41023 112289 41051
rect 112323 41023 112351 41051
rect 112137 40961 112165 40989
rect 112199 40961 112227 40989
rect 112261 40961 112289 40989
rect 112323 40961 112351 40989
rect 112137 32147 112165 32175
rect 112199 32147 112227 32175
rect 112261 32147 112289 32175
rect 112323 32147 112351 32175
rect 112137 32085 112165 32113
rect 112199 32085 112227 32113
rect 112261 32085 112289 32113
rect 112323 32085 112351 32113
rect 112137 32023 112165 32051
rect 112199 32023 112227 32051
rect 112261 32023 112289 32051
rect 112323 32023 112351 32051
rect 112137 31961 112165 31989
rect 112199 31961 112227 31989
rect 112261 31961 112289 31989
rect 112323 31961 112351 31989
rect 112137 23147 112165 23175
rect 112199 23147 112227 23175
rect 112261 23147 112289 23175
rect 112323 23147 112351 23175
rect 112137 23085 112165 23113
rect 112199 23085 112227 23113
rect 112261 23085 112289 23113
rect 112323 23085 112351 23113
rect 112137 23023 112165 23051
rect 112199 23023 112227 23051
rect 112261 23023 112289 23051
rect 112323 23023 112351 23051
rect 112137 22961 112165 22989
rect 112199 22961 112227 22989
rect 112261 22961 112289 22989
rect 112323 22961 112351 22989
rect 112137 14147 112165 14175
rect 112199 14147 112227 14175
rect 112261 14147 112289 14175
rect 112323 14147 112351 14175
rect 112137 14085 112165 14113
rect 112199 14085 112227 14113
rect 112261 14085 112289 14113
rect 112323 14085 112351 14113
rect 112137 14023 112165 14051
rect 112199 14023 112227 14051
rect 112261 14023 112289 14051
rect 112323 14023 112351 14051
rect 112137 13961 112165 13989
rect 112199 13961 112227 13989
rect 112261 13961 112289 13989
rect 112323 13961 112351 13989
rect 112137 5147 112165 5175
rect 112199 5147 112227 5175
rect 112261 5147 112289 5175
rect 112323 5147 112351 5175
rect 112137 5085 112165 5113
rect 112199 5085 112227 5113
rect 112261 5085 112289 5113
rect 112323 5085 112351 5113
rect 112137 5023 112165 5051
rect 112199 5023 112227 5051
rect 112261 5023 112289 5051
rect 112323 5023 112351 5051
rect 112137 4961 112165 4989
rect 112199 4961 112227 4989
rect 112261 4961 112289 4989
rect 112323 4961 112351 4989
rect 112137 -588 112165 -560
rect 112199 -588 112227 -560
rect 112261 -588 112289 -560
rect 112323 -588 112351 -560
rect 112137 -650 112165 -622
rect 112199 -650 112227 -622
rect 112261 -650 112289 -622
rect 112323 -650 112351 -622
rect 112137 -712 112165 -684
rect 112199 -712 112227 -684
rect 112261 -712 112289 -684
rect 112323 -712 112351 -684
rect 112137 -774 112165 -746
rect 112199 -774 112227 -746
rect 112261 -774 112289 -746
rect 112323 -774 112351 -746
rect 125637 92147 125665 92175
rect 125699 92147 125727 92175
rect 125761 92147 125789 92175
rect 125823 92147 125851 92175
rect 125637 92085 125665 92113
rect 125699 92085 125727 92113
rect 125761 92085 125789 92113
rect 125823 92085 125851 92113
rect 125637 92023 125665 92051
rect 125699 92023 125727 92051
rect 125761 92023 125789 92051
rect 125823 92023 125851 92051
rect 125637 91961 125665 91989
rect 125699 91961 125727 91989
rect 125761 91961 125789 91989
rect 125823 91961 125851 91989
rect 125637 83147 125665 83175
rect 125699 83147 125727 83175
rect 125761 83147 125789 83175
rect 125823 83147 125851 83175
rect 125637 83085 125665 83113
rect 125699 83085 125727 83113
rect 125761 83085 125789 83113
rect 125823 83085 125851 83113
rect 125637 83023 125665 83051
rect 125699 83023 125727 83051
rect 125761 83023 125789 83051
rect 125823 83023 125851 83051
rect 125637 82961 125665 82989
rect 125699 82961 125727 82989
rect 125761 82961 125789 82989
rect 125823 82961 125851 82989
rect 125637 74147 125665 74175
rect 125699 74147 125727 74175
rect 125761 74147 125789 74175
rect 125823 74147 125851 74175
rect 125637 74085 125665 74113
rect 125699 74085 125727 74113
rect 125761 74085 125789 74113
rect 125823 74085 125851 74113
rect 125637 74023 125665 74051
rect 125699 74023 125727 74051
rect 125761 74023 125789 74051
rect 125823 74023 125851 74051
rect 125637 73961 125665 73989
rect 125699 73961 125727 73989
rect 125761 73961 125789 73989
rect 125823 73961 125851 73989
rect 125637 65147 125665 65175
rect 125699 65147 125727 65175
rect 125761 65147 125789 65175
rect 125823 65147 125851 65175
rect 125637 65085 125665 65113
rect 125699 65085 125727 65113
rect 125761 65085 125789 65113
rect 125823 65085 125851 65113
rect 125637 65023 125665 65051
rect 125699 65023 125727 65051
rect 125761 65023 125789 65051
rect 125823 65023 125851 65051
rect 125637 64961 125665 64989
rect 125699 64961 125727 64989
rect 125761 64961 125789 64989
rect 125823 64961 125851 64989
rect 125637 56147 125665 56175
rect 125699 56147 125727 56175
rect 125761 56147 125789 56175
rect 125823 56147 125851 56175
rect 125637 56085 125665 56113
rect 125699 56085 125727 56113
rect 125761 56085 125789 56113
rect 125823 56085 125851 56113
rect 125637 56023 125665 56051
rect 125699 56023 125727 56051
rect 125761 56023 125789 56051
rect 125823 56023 125851 56051
rect 125637 55961 125665 55989
rect 125699 55961 125727 55989
rect 125761 55961 125789 55989
rect 125823 55961 125851 55989
rect 125637 47147 125665 47175
rect 125699 47147 125727 47175
rect 125761 47147 125789 47175
rect 125823 47147 125851 47175
rect 125637 47085 125665 47113
rect 125699 47085 125727 47113
rect 125761 47085 125789 47113
rect 125823 47085 125851 47113
rect 125637 47023 125665 47051
rect 125699 47023 125727 47051
rect 125761 47023 125789 47051
rect 125823 47023 125851 47051
rect 125637 46961 125665 46989
rect 125699 46961 125727 46989
rect 125761 46961 125789 46989
rect 125823 46961 125851 46989
rect 125637 38147 125665 38175
rect 125699 38147 125727 38175
rect 125761 38147 125789 38175
rect 125823 38147 125851 38175
rect 125637 38085 125665 38113
rect 125699 38085 125727 38113
rect 125761 38085 125789 38113
rect 125823 38085 125851 38113
rect 125637 38023 125665 38051
rect 125699 38023 125727 38051
rect 125761 38023 125789 38051
rect 125823 38023 125851 38051
rect 125637 37961 125665 37989
rect 125699 37961 125727 37989
rect 125761 37961 125789 37989
rect 125823 37961 125851 37989
rect 125637 29147 125665 29175
rect 125699 29147 125727 29175
rect 125761 29147 125789 29175
rect 125823 29147 125851 29175
rect 125637 29085 125665 29113
rect 125699 29085 125727 29113
rect 125761 29085 125789 29113
rect 125823 29085 125851 29113
rect 125637 29023 125665 29051
rect 125699 29023 125727 29051
rect 125761 29023 125789 29051
rect 125823 29023 125851 29051
rect 125637 28961 125665 28989
rect 125699 28961 125727 28989
rect 125761 28961 125789 28989
rect 125823 28961 125851 28989
rect 125637 20147 125665 20175
rect 125699 20147 125727 20175
rect 125761 20147 125789 20175
rect 125823 20147 125851 20175
rect 125637 20085 125665 20113
rect 125699 20085 125727 20113
rect 125761 20085 125789 20113
rect 125823 20085 125851 20113
rect 125637 20023 125665 20051
rect 125699 20023 125727 20051
rect 125761 20023 125789 20051
rect 125823 20023 125851 20051
rect 125637 19961 125665 19989
rect 125699 19961 125727 19989
rect 125761 19961 125789 19989
rect 125823 19961 125851 19989
rect 125637 11147 125665 11175
rect 125699 11147 125727 11175
rect 125761 11147 125789 11175
rect 125823 11147 125851 11175
rect 125637 11085 125665 11113
rect 125699 11085 125727 11113
rect 125761 11085 125789 11113
rect 125823 11085 125851 11113
rect 125637 11023 125665 11051
rect 125699 11023 125727 11051
rect 125761 11023 125789 11051
rect 125823 11023 125851 11051
rect 125637 10961 125665 10989
rect 125699 10961 125727 10989
rect 125761 10961 125789 10989
rect 125823 10961 125851 10989
rect 125637 2147 125665 2175
rect 125699 2147 125727 2175
rect 125761 2147 125789 2175
rect 125823 2147 125851 2175
rect 125637 2085 125665 2113
rect 125699 2085 125727 2113
rect 125761 2085 125789 2113
rect 125823 2085 125851 2113
rect 125637 2023 125665 2051
rect 125699 2023 125727 2051
rect 125761 2023 125789 2051
rect 125823 2023 125851 2051
rect 125637 1961 125665 1989
rect 125699 1961 125727 1989
rect 125761 1961 125789 1989
rect 125823 1961 125851 1989
rect 125637 -108 125665 -80
rect 125699 -108 125727 -80
rect 125761 -108 125789 -80
rect 125823 -108 125851 -80
rect 125637 -170 125665 -142
rect 125699 -170 125727 -142
rect 125761 -170 125789 -142
rect 125823 -170 125851 -142
rect 125637 -232 125665 -204
rect 125699 -232 125727 -204
rect 125761 -232 125789 -204
rect 125823 -232 125851 -204
rect 125637 -294 125665 -266
rect 125699 -294 125727 -266
rect 125761 -294 125789 -266
rect 125823 -294 125851 -266
rect 127497 130986 127525 131014
rect 127559 130986 127587 131014
rect 127621 130986 127649 131014
rect 127683 130986 127711 131014
rect 127497 130924 127525 130952
rect 127559 130924 127587 130952
rect 127621 130924 127649 130952
rect 127683 130924 127711 130952
rect 127497 122147 127525 122175
rect 127559 122147 127587 122175
rect 127621 122147 127649 122175
rect 127683 122147 127711 122175
rect 127497 122085 127525 122113
rect 127559 122085 127587 122113
rect 127621 122085 127649 122113
rect 127683 122085 127711 122113
rect 127497 122023 127525 122051
rect 127559 122023 127587 122051
rect 127621 122023 127649 122051
rect 127683 122023 127711 122051
rect 127497 121961 127525 121989
rect 127559 121961 127587 121989
rect 127621 121961 127649 121989
rect 127683 121961 127711 121989
rect 127497 113147 127525 113175
rect 127559 113147 127587 113175
rect 127621 113147 127649 113175
rect 127683 113147 127711 113175
rect 127497 113085 127525 113113
rect 127559 113085 127587 113113
rect 127621 113085 127649 113113
rect 127683 113085 127711 113113
rect 127497 113023 127525 113051
rect 127559 113023 127587 113051
rect 127621 113023 127649 113051
rect 127683 113023 127711 113051
rect 127497 112961 127525 112989
rect 127559 112961 127587 112989
rect 127621 112961 127649 112989
rect 127683 112961 127711 112989
rect 127497 104147 127525 104175
rect 127559 104147 127587 104175
rect 127621 104147 127649 104175
rect 127683 104147 127711 104175
rect 127497 104085 127525 104113
rect 127559 104085 127587 104113
rect 127621 104085 127649 104113
rect 127683 104085 127711 104113
rect 127497 104023 127525 104051
rect 127559 104023 127587 104051
rect 127621 104023 127649 104051
rect 127683 104023 127711 104051
rect 127497 103961 127525 103989
rect 127559 103961 127587 103989
rect 127621 103961 127649 103989
rect 127683 103961 127711 103989
rect 127497 95147 127525 95175
rect 127559 95147 127587 95175
rect 127621 95147 127649 95175
rect 127683 95147 127711 95175
rect 127497 95085 127525 95113
rect 127559 95085 127587 95113
rect 127621 95085 127649 95113
rect 127683 95085 127711 95113
rect 127497 95023 127525 95051
rect 127559 95023 127587 95051
rect 127621 95023 127649 95051
rect 127683 95023 127711 95051
rect 127497 94961 127525 94989
rect 127559 94961 127587 94989
rect 127621 94961 127649 94989
rect 127683 94961 127711 94989
rect 127497 86147 127525 86175
rect 127559 86147 127587 86175
rect 127621 86147 127649 86175
rect 127683 86147 127711 86175
rect 127497 86085 127525 86113
rect 127559 86085 127587 86113
rect 127621 86085 127649 86113
rect 127683 86085 127711 86113
rect 127497 86023 127525 86051
rect 127559 86023 127587 86051
rect 127621 86023 127649 86051
rect 127683 86023 127711 86051
rect 127497 85961 127525 85989
rect 127559 85961 127587 85989
rect 127621 85961 127649 85989
rect 127683 85961 127711 85989
rect 127497 77147 127525 77175
rect 127559 77147 127587 77175
rect 127621 77147 127649 77175
rect 127683 77147 127711 77175
rect 127497 77085 127525 77113
rect 127559 77085 127587 77113
rect 127621 77085 127649 77113
rect 127683 77085 127711 77113
rect 127497 77023 127525 77051
rect 127559 77023 127587 77051
rect 127621 77023 127649 77051
rect 127683 77023 127711 77051
rect 127497 76961 127525 76989
rect 127559 76961 127587 76989
rect 127621 76961 127649 76989
rect 127683 76961 127711 76989
rect 127497 68147 127525 68175
rect 127559 68147 127587 68175
rect 127621 68147 127649 68175
rect 127683 68147 127711 68175
rect 127497 68085 127525 68113
rect 127559 68085 127587 68113
rect 127621 68085 127649 68113
rect 127683 68085 127711 68113
rect 127497 68023 127525 68051
rect 127559 68023 127587 68051
rect 127621 68023 127649 68051
rect 127683 68023 127711 68051
rect 127497 67961 127525 67989
rect 127559 67961 127587 67989
rect 127621 67961 127649 67989
rect 127683 67961 127711 67989
rect 127497 59147 127525 59175
rect 127559 59147 127587 59175
rect 127621 59147 127649 59175
rect 127683 59147 127711 59175
rect 127497 59085 127525 59113
rect 127559 59085 127587 59113
rect 127621 59085 127649 59113
rect 127683 59085 127711 59113
rect 127497 59023 127525 59051
rect 127559 59023 127587 59051
rect 127621 59023 127649 59051
rect 127683 59023 127711 59051
rect 127497 58961 127525 58989
rect 127559 58961 127587 58989
rect 127621 58961 127649 58989
rect 127683 58961 127711 58989
rect 127497 50147 127525 50175
rect 127559 50147 127587 50175
rect 127621 50147 127649 50175
rect 127683 50147 127711 50175
rect 127497 50085 127525 50113
rect 127559 50085 127587 50113
rect 127621 50085 127649 50113
rect 127683 50085 127711 50113
rect 127497 50023 127525 50051
rect 127559 50023 127587 50051
rect 127621 50023 127649 50051
rect 127683 50023 127711 50051
rect 127497 49961 127525 49989
rect 127559 49961 127587 49989
rect 127621 49961 127649 49989
rect 127683 49961 127711 49989
rect 127497 41147 127525 41175
rect 127559 41147 127587 41175
rect 127621 41147 127649 41175
rect 127683 41147 127711 41175
rect 127497 41085 127525 41113
rect 127559 41085 127587 41113
rect 127621 41085 127649 41113
rect 127683 41085 127711 41113
rect 127497 41023 127525 41051
rect 127559 41023 127587 41051
rect 127621 41023 127649 41051
rect 127683 41023 127711 41051
rect 127497 40961 127525 40989
rect 127559 40961 127587 40989
rect 127621 40961 127649 40989
rect 127683 40961 127711 40989
rect 127497 32147 127525 32175
rect 127559 32147 127587 32175
rect 127621 32147 127649 32175
rect 127683 32147 127711 32175
rect 127497 32085 127525 32113
rect 127559 32085 127587 32113
rect 127621 32085 127649 32113
rect 127683 32085 127711 32113
rect 127497 32023 127525 32051
rect 127559 32023 127587 32051
rect 127621 32023 127649 32051
rect 127683 32023 127711 32051
rect 127497 31961 127525 31989
rect 127559 31961 127587 31989
rect 127621 31961 127649 31989
rect 127683 31961 127711 31989
rect 127497 23147 127525 23175
rect 127559 23147 127587 23175
rect 127621 23147 127649 23175
rect 127683 23147 127711 23175
rect 127497 23085 127525 23113
rect 127559 23085 127587 23113
rect 127621 23085 127649 23113
rect 127683 23085 127711 23113
rect 127497 23023 127525 23051
rect 127559 23023 127587 23051
rect 127621 23023 127649 23051
rect 127683 23023 127711 23051
rect 127497 22961 127525 22989
rect 127559 22961 127587 22989
rect 127621 22961 127649 22989
rect 127683 22961 127711 22989
rect 127497 14147 127525 14175
rect 127559 14147 127587 14175
rect 127621 14147 127649 14175
rect 127683 14147 127711 14175
rect 127497 14085 127525 14113
rect 127559 14085 127587 14113
rect 127621 14085 127649 14113
rect 127683 14085 127711 14113
rect 127497 14023 127525 14051
rect 127559 14023 127587 14051
rect 127621 14023 127649 14051
rect 127683 14023 127711 14051
rect 127497 13961 127525 13989
rect 127559 13961 127587 13989
rect 127621 13961 127649 13989
rect 127683 13961 127711 13989
rect 127497 5147 127525 5175
rect 127559 5147 127587 5175
rect 127621 5147 127649 5175
rect 127683 5147 127711 5175
rect 127497 5085 127525 5113
rect 127559 5085 127587 5113
rect 127621 5085 127649 5113
rect 127683 5085 127711 5113
rect 127497 5023 127525 5051
rect 127559 5023 127587 5051
rect 127621 5023 127649 5051
rect 127683 5023 127711 5051
rect 127497 4961 127525 4989
rect 127559 4961 127587 4989
rect 127621 4961 127649 4989
rect 127683 4961 127711 4989
rect 127497 -588 127525 -560
rect 127559 -588 127587 -560
rect 127621 -588 127649 -560
rect 127683 -588 127711 -560
rect 127497 -650 127525 -622
rect 127559 -650 127587 -622
rect 127621 -650 127649 -622
rect 127683 -650 127711 -622
rect 127497 -712 127525 -684
rect 127559 -712 127587 -684
rect 127621 -712 127649 -684
rect 127683 -712 127711 -684
rect 127497 -774 127525 -746
rect 127559 -774 127587 -746
rect 127621 -774 127649 -746
rect 127683 -774 127711 -746
rect 140997 128147 141025 128175
rect 141059 128147 141087 128175
rect 141121 128147 141149 128175
rect 141183 128147 141211 128175
rect 140997 128085 141025 128113
rect 141059 128085 141087 128113
rect 141121 128085 141149 128113
rect 141183 128085 141211 128113
rect 140997 128023 141025 128051
rect 141059 128023 141087 128051
rect 141121 128023 141149 128051
rect 141183 128023 141211 128051
rect 140997 127961 141025 127989
rect 141059 127961 141087 127989
rect 141121 127961 141149 127989
rect 141183 127961 141211 127989
rect 140997 119147 141025 119175
rect 141059 119147 141087 119175
rect 141121 119147 141149 119175
rect 141183 119147 141211 119175
rect 140997 119085 141025 119113
rect 141059 119085 141087 119113
rect 141121 119085 141149 119113
rect 141183 119085 141211 119113
rect 140997 119023 141025 119051
rect 141059 119023 141087 119051
rect 141121 119023 141149 119051
rect 141183 119023 141211 119051
rect 140997 118961 141025 118989
rect 141059 118961 141087 118989
rect 141121 118961 141149 118989
rect 141183 118961 141211 118989
rect 140997 110147 141025 110175
rect 141059 110147 141087 110175
rect 141121 110147 141149 110175
rect 141183 110147 141211 110175
rect 140997 110085 141025 110113
rect 141059 110085 141087 110113
rect 141121 110085 141149 110113
rect 141183 110085 141211 110113
rect 140997 110023 141025 110051
rect 141059 110023 141087 110051
rect 141121 110023 141149 110051
rect 141183 110023 141211 110051
rect 140997 109961 141025 109989
rect 141059 109961 141087 109989
rect 141121 109961 141149 109989
rect 141183 109961 141211 109989
rect 140997 101147 141025 101175
rect 141059 101147 141087 101175
rect 141121 101147 141149 101175
rect 141183 101147 141211 101175
rect 140997 101085 141025 101113
rect 141059 101085 141087 101113
rect 141121 101085 141149 101113
rect 141183 101085 141211 101113
rect 140997 101023 141025 101051
rect 141059 101023 141087 101051
rect 141121 101023 141149 101051
rect 141183 101023 141211 101051
rect 140997 100961 141025 100989
rect 141059 100961 141087 100989
rect 141121 100961 141149 100989
rect 141183 100961 141211 100989
rect 140997 92147 141025 92175
rect 141059 92147 141087 92175
rect 141121 92147 141149 92175
rect 141183 92147 141211 92175
rect 140997 92085 141025 92113
rect 141059 92085 141087 92113
rect 141121 92085 141149 92113
rect 141183 92085 141211 92113
rect 140997 92023 141025 92051
rect 141059 92023 141087 92051
rect 141121 92023 141149 92051
rect 141183 92023 141211 92051
rect 140997 91961 141025 91989
rect 141059 91961 141087 91989
rect 141121 91961 141149 91989
rect 141183 91961 141211 91989
rect 140997 83147 141025 83175
rect 141059 83147 141087 83175
rect 141121 83147 141149 83175
rect 141183 83147 141211 83175
rect 140997 83085 141025 83113
rect 141059 83085 141087 83113
rect 141121 83085 141149 83113
rect 141183 83085 141211 83113
rect 140997 83023 141025 83051
rect 141059 83023 141087 83051
rect 141121 83023 141149 83051
rect 141183 83023 141211 83051
rect 140997 82961 141025 82989
rect 141059 82961 141087 82989
rect 141121 82961 141149 82989
rect 141183 82961 141211 82989
rect 140997 74147 141025 74175
rect 141059 74147 141087 74175
rect 141121 74147 141149 74175
rect 141183 74147 141211 74175
rect 140997 74085 141025 74113
rect 141059 74085 141087 74113
rect 141121 74085 141149 74113
rect 141183 74085 141211 74113
rect 140997 74023 141025 74051
rect 141059 74023 141087 74051
rect 141121 74023 141149 74051
rect 141183 74023 141211 74051
rect 140997 73961 141025 73989
rect 141059 73961 141087 73989
rect 141121 73961 141149 73989
rect 141183 73961 141211 73989
rect 140997 65147 141025 65175
rect 141059 65147 141087 65175
rect 141121 65147 141149 65175
rect 141183 65147 141211 65175
rect 140997 65085 141025 65113
rect 141059 65085 141087 65113
rect 141121 65085 141149 65113
rect 141183 65085 141211 65113
rect 140997 65023 141025 65051
rect 141059 65023 141087 65051
rect 141121 65023 141149 65051
rect 141183 65023 141211 65051
rect 140997 64961 141025 64989
rect 141059 64961 141087 64989
rect 141121 64961 141149 64989
rect 141183 64961 141211 64989
rect 140997 56147 141025 56175
rect 141059 56147 141087 56175
rect 141121 56147 141149 56175
rect 141183 56147 141211 56175
rect 140997 56085 141025 56113
rect 141059 56085 141087 56113
rect 141121 56085 141149 56113
rect 141183 56085 141211 56113
rect 140997 56023 141025 56051
rect 141059 56023 141087 56051
rect 141121 56023 141149 56051
rect 141183 56023 141211 56051
rect 140997 55961 141025 55989
rect 141059 55961 141087 55989
rect 141121 55961 141149 55989
rect 141183 55961 141211 55989
rect 140997 47147 141025 47175
rect 141059 47147 141087 47175
rect 141121 47147 141149 47175
rect 141183 47147 141211 47175
rect 140997 47085 141025 47113
rect 141059 47085 141087 47113
rect 141121 47085 141149 47113
rect 141183 47085 141211 47113
rect 140997 47023 141025 47051
rect 141059 47023 141087 47051
rect 141121 47023 141149 47051
rect 141183 47023 141211 47051
rect 140997 46961 141025 46989
rect 141059 46961 141087 46989
rect 141121 46961 141149 46989
rect 141183 46961 141211 46989
rect 140997 38147 141025 38175
rect 141059 38147 141087 38175
rect 141121 38147 141149 38175
rect 141183 38147 141211 38175
rect 140997 38085 141025 38113
rect 141059 38085 141087 38113
rect 141121 38085 141149 38113
rect 141183 38085 141211 38113
rect 140997 38023 141025 38051
rect 141059 38023 141087 38051
rect 141121 38023 141149 38051
rect 141183 38023 141211 38051
rect 140997 37961 141025 37989
rect 141059 37961 141087 37989
rect 141121 37961 141149 37989
rect 141183 37961 141211 37989
rect 140997 29147 141025 29175
rect 141059 29147 141087 29175
rect 141121 29147 141149 29175
rect 141183 29147 141211 29175
rect 140997 29085 141025 29113
rect 141059 29085 141087 29113
rect 141121 29085 141149 29113
rect 141183 29085 141211 29113
rect 140997 29023 141025 29051
rect 141059 29023 141087 29051
rect 141121 29023 141149 29051
rect 141183 29023 141211 29051
rect 140997 28961 141025 28989
rect 141059 28961 141087 28989
rect 141121 28961 141149 28989
rect 141183 28961 141211 28989
rect 140997 20147 141025 20175
rect 141059 20147 141087 20175
rect 141121 20147 141149 20175
rect 141183 20147 141211 20175
rect 140997 20085 141025 20113
rect 141059 20085 141087 20113
rect 141121 20085 141149 20113
rect 141183 20085 141211 20113
rect 140997 20023 141025 20051
rect 141059 20023 141087 20051
rect 141121 20023 141149 20051
rect 141183 20023 141211 20051
rect 140997 19961 141025 19989
rect 141059 19961 141087 19989
rect 141121 19961 141149 19989
rect 141183 19961 141211 19989
rect 140997 11147 141025 11175
rect 141059 11147 141087 11175
rect 141121 11147 141149 11175
rect 141183 11147 141211 11175
rect 140997 11085 141025 11113
rect 141059 11085 141087 11113
rect 141121 11085 141149 11113
rect 141183 11085 141211 11113
rect 140997 11023 141025 11051
rect 141059 11023 141087 11051
rect 141121 11023 141149 11051
rect 141183 11023 141211 11051
rect 140997 10961 141025 10989
rect 141059 10961 141087 10989
rect 141121 10961 141149 10989
rect 141183 10961 141211 10989
rect 140997 2147 141025 2175
rect 141059 2147 141087 2175
rect 141121 2147 141149 2175
rect 141183 2147 141211 2175
rect 140997 2085 141025 2113
rect 141059 2085 141087 2113
rect 141121 2085 141149 2113
rect 141183 2085 141211 2113
rect 140997 2023 141025 2051
rect 141059 2023 141087 2051
rect 141121 2023 141149 2051
rect 141183 2023 141211 2051
rect 140997 1961 141025 1989
rect 141059 1961 141087 1989
rect 141121 1961 141149 1989
rect 141183 1961 141211 1989
rect 140997 -108 141025 -80
rect 141059 -108 141087 -80
rect 141121 -108 141149 -80
rect 141183 -108 141211 -80
rect 140997 -170 141025 -142
rect 141059 -170 141087 -142
rect 141121 -170 141149 -142
rect 141183 -170 141211 -142
rect 140997 -232 141025 -204
rect 141059 -232 141087 -204
rect 141121 -232 141149 -204
rect 141183 -232 141211 -204
rect 140997 -294 141025 -266
rect 141059 -294 141087 -266
rect 141121 -294 141149 -266
rect 141183 -294 141211 -266
rect 142857 130986 142885 131014
rect 142919 130986 142947 131014
rect 142981 130986 143009 131014
rect 143043 130986 143071 131014
rect 142857 130924 142885 130952
rect 142919 130924 142947 130952
rect 142981 130924 143009 130952
rect 143043 130924 143071 130952
rect 142857 122147 142885 122175
rect 142919 122147 142947 122175
rect 142981 122147 143009 122175
rect 143043 122147 143071 122175
rect 142857 122085 142885 122113
rect 142919 122085 142947 122113
rect 142981 122085 143009 122113
rect 143043 122085 143071 122113
rect 142857 122023 142885 122051
rect 142919 122023 142947 122051
rect 142981 122023 143009 122051
rect 143043 122023 143071 122051
rect 142857 121961 142885 121989
rect 142919 121961 142947 121989
rect 142981 121961 143009 121989
rect 143043 121961 143071 121989
rect 142857 113147 142885 113175
rect 142919 113147 142947 113175
rect 142981 113147 143009 113175
rect 143043 113147 143071 113175
rect 142857 113085 142885 113113
rect 142919 113085 142947 113113
rect 142981 113085 143009 113113
rect 143043 113085 143071 113113
rect 142857 113023 142885 113051
rect 142919 113023 142947 113051
rect 142981 113023 143009 113051
rect 143043 113023 143071 113051
rect 142857 112961 142885 112989
rect 142919 112961 142947 112989
rect 142981 112961 143009 112989
rect 143043 112961 143071 112989
rect 142857 104147 142885 104175
rect 142919 104147 142947 104175
rect 142981 104147 143009 104175
rect 143043 104147 143071 104175
rect 142857 104085 142885 104113
rect 142919 104085 142947 104113
rect 142981 104085 143009 104113
rect 143043 104085 143071 104113
rect 142857 104023 142885 104051
rect 142919 104023 142947 104051
rect 142981 104023 143009 104051
rect 143043 104023 143071 104051
rect 142857 103961 142885 103989
rect 142919 103961 142947 103989
rect 142981 103961 143009 103989
rect 143043 103961 143071 103989
rect 142857 95147 142885 95175
rect 142919 95147 142947 95175
rect 142981 95147 143009 95175
rect 143043 95147 143071 95175
rect 142857 95085 142885 95113
rect 142919 95085 142947 95113
rect 142981 95085 143009 95113
rect 143043 95085 143071 95113
rect 142857 95023 142885 95051
rect 142919 95023 142947 95051
rect 142981 95023 143009 95051
rect 143043 95023 143071 95051
rect 142857 94961 142885 94989
rect 142919 94961 142947 94989
rect 142981 94961 143009 94989
rect 143043 94961 143071 94989
rect 142857 86147 142885 86175
rect 142919 86147 142947 86175
rect 142981 86147 143009 86175
rect 143043 86147 143071 86175
rect 142857 86085 142885 86113
rect 142919 86085 142947 86113
rect 142981 86085 143009 86113
rect 143043 86085 143071 86113
rect 142857 86023 142885 86051
rect 142919 86023 142947 86051
rect 142981 86023 143009 86051
rect 143043 86023 143071 86051
rect 142857 85961 142885 85989
rect 142919 85961 142947 85989
rect 142981 85961 143009 85989
rect 143043 85961 143071 85989
rect 142857 77147 142885 77175
rect 142919 77147 142947 77175
rect 142981 77147 143009 77175
rect 143043 77147 143071 77175
rect 142857 77085 142885 77113
rect 142919 77085 142947 77113
rect 142981 77085 143009 77113
rect 143043 77085 143071 77113
rect 142857 77023 142885 77051
rect 142919 77023 142947 77051
rect 142981 77023 143009 77051
rect 143043 77023 143071 77051
rect 142857 76961 142885 76989
rect 142919 76961 142947 76989
rect 142981 76961 143009 76989
rect 143043 76961 143071 76989
rect 142857 68147 142885 68175
rect 142919 68147 142947 68175
rect 142981 68147 143009 68175
rect 143043 68147 143071 68175
rect 142857 68085 142885 68113
rect 142919 68085 142947 68113
rect 142981 68085 143009 68113
rect 143043 68085 143071 68113
rect 142857 68023 142885 68051
rect 142919 68023 142947 68051
rect 142981 68023 143009 68051
rect 143043 68023 143071 68051
rect 142857 67961 142885 67989
rect 142919 67961 142947 67989
rect 142981 67961 143009 67989
rect 143043 67961 143071 67989
rect 142857 59147 142885 59175
rect 142919 59147 142947 59175
rect 142981 59147 143009 59175
rect 143043 59147 143071 59175
rect 142857 59085 142885 59113
rect 142919 59085 142947 59113
rect 142981 59085 143009 59113
rect 143043 59085 143071 59113
rect 142857 59023 142885 59051
rect 142919 59023 142947 59051
rect 142981 59023 143009 59051
rect 143043 59023 143071 59051
rect 142857 58961 142885 58989
rect 142919 58961 142947 58989
rect 142981 58961 143009 58989
rect 143043 58961 143071 58989
rect 142857 50147 142885 50175
rect 142919 50147 142947 50175
rect 142981 50147 143009 50175
rect 143043 50147 143071 50175
rect 142857 50085 142885 50113
rect 142919 50085 142947 50113
rect 142981 50085 143009 50113
rect 143043 50085 143071 50113
rect 142857 50023 142885 50051
rect 142919 50023 142947 50051
rect 142981 50023 143009 50051
rect 143043 50023 143071 50051
rect 142857 49961 142885 49989
rect 142919 49961 142947 49989
rect 142981 49961 143009 49989
rect 143043 49961 143071 49989
rect 142857 41147 142885 41175
rect 142919 41147 142947 41175
rect 142981 41147 143009 41175
rect 143043 41147 143071 41175
rect 142857 41085 142885 41113
rect 142919 41085 142947 41113
rect 142981 41085 143009 41113
rect 143043 41085 143071 41113
rect 142857 41023 142885 41051
rect 142919 41023 142947 41051
rect 142981 41023 143009 41051
rect 143043 41023 143071 41051
rect 142857 40961 142885 40989
rect 142919 40961 142947 40989
rect 142981 40961 143009 40989
rect 143043 40961 143071 40989
rect 142857 32147 142885 32175
rect 142919 32147 142947 32175
rect 142981 32147 143009 32175
rect 143043 32147 143071 32175
rect 142857 32085 142885 32113
rect 142919 32085 142947 32113
rect 142981 32085 143009 32113
rect 143043 32085 143071 32113
rect 142857 32023 142885 32051
rect 142919 32023 142947 32051
rect 142981 32023 143009 32051
rect 143043 32023 143071 32051
rect 142857 31961 142885 31989
rect 142919 31961 142947 31989
rect 142981 31961 143009 31989
rect 143043 31961 143071 31989
rect 142857 23147 142885 23175
rect 142919 23147 142947 23175
rect 142981 23147 143009 23175
rect 143043 23147 143071 23175
rect 142857 23085 142885 23113
rect 142919 23085 142947 23113
rect 142981 23085 143009 23113
rect 143043 23085 143071 23113
rect 142857 23023 142885 23051
rect 142919 23023 142947 23051
rect 142981 23023 143009 23051
rect 143043 23023 143071 23051
rect 142857 22961 142885 22989
rect 142919 22961 142947 22989
rect 142981 22961 143009 22989
rect 143043 22961 143071 22989
rect 142857 14147 142885 14175
rect 142919 14147 142947 14175
rect 142981 14147 143009 14175
rect 143043 14147 143071 14175
rect 142857 14085 142885 14113
rect 142919 14085 142947 14113
rect 142981 14085 143009 14113
rect 143043 14085 143071 14113
rect 142857 14023 142885 14051
rect 142919 14023 142947 14051
rect 142981 14023 143009 14051
rect 143043 14023 143071 14051
rect 142857 13961 142885 13989
rect 142919 13961 142947 13989
rect 142981 13961 143009 13989
rect 143043 13961 143071 13989
rect 142857 5147 142885 5175
rect 142919 5147 142947 5175
rect 142981 5147 143009 5175
rect 143043 5147 143071 5175
rect 142857 5085 142885 5113
rect 142919 5085 142947 5113
rect 142981 5085 143009 5113
rect 143043 5085 143071 5113
rect 142857 5023 142885 5051
rect 142919 5023 142947 5051
rect 142981 5023 143009 5051
rect 143043 5023 143071 5051
rect 142857 4961 142885 4989
rect 142919 4961 142947 4989
rect 142981 4961 143009 4989
rect 143043 4961 143071 4989
rect 142857 -588 142885 -560
rect 142919 -588 142947 -560
rect 142981 -588 143009 -560
rect 143043 -588 143071 -560
rect 142857 -650 142885 -622
rect 142919 -650 142947 -622
rect 142981 -650 143009 -622
rect 143043 -650 143071 -622
rect 142857 -712 142885 -684
rect 142919 -712 142947 -684
rect 142981 -712 143009 -684
rect 143043 -712 143071 -684
rect 142857 -774 142885 -746
rect 142919 -774 142947 -746
rect 142981 -774 143009 -746
rect 143043 -774 143071 -746
rect 156357 128147 156385 128175
rect 156419 128147 156447 128175
rect 156481 128147 156509 128175
rect 156543 128147 156571 128175
rect 156357 128085 156385 128113
rect 156419 128085 156447 128113
rect 156481 128085 156509 128113
rect 156543 128085 156571 128113
rect 156357 128023 156385 128051
rect 156419 128023 156447 128051
rect 156481 128023 156509 128051
rect 156543 128023 156571 128051
rect 156357 127961 156385 127989
rect 156419 127961 156447 127989
rect 156481 127961 156509 127989
rect 156543 127961 156571 127989
rect 156357 119147 156385 119175
rect 156419 119147 156447 119175
rect 156481 119147 156509 119175
rect 156543 119147 156571 119175
rect 156357 119085 156385 119113
rect 156419 119085 156447 119113
rect 156481 119085 156509 119113
rect 156543 119085 156571 119113
rect 156357 119023 156385 119051
rect 156419 119023 156447 119051
rect 156481 119023 156509 119051
rect 156543 119023 156571 119051
rect 156357 118961 156385 118989
rect 156419 118961 156447 118989
rect 156481 118961 156509 118989
rect 156543 118961 156571 118989
rect 156357 110147 156385 110175
rect 156419 110147 156447 110175
rect 156481 110147 156509 110175
rect 156543 110147 156571 110175
rect 156357 110085 156385 110113
rect 156419 110085 156447 110113
rect 156481 110085 156509 110113
rect 156543 110085 156571 110113
rect 156357 110023 156385 110051
rect 156419 110023 156447 110051
rect 156481 110023 156509 110051
rect 156543 110023 156571 110051
rect 156357 109961 156385 109989
rect 156419 109961 156447 109989
rect 156481 109961 156509 109989
rect 156543 109961 156571 109989
rect 156357 101147 156385 101175
rect 156419 101147 156447 101175
rect 156481 101147 156509 101175
rect 156543 101147 156571 101175
rect 156357 101085 156385 101113
rect 156419 101085 156447 101113
rect 156481 101085 156509 101113
rect 156543 101085 156571 101113
rect 156357 101023 156385 101051
rect 156419 101023 156447 101051
rect 156481 101023 156509 101051
rect 156543 101023 156571 101051
rect 156357 100961 156385 100989
rect 156419 100961 156447 100989
rect 156481 100961 156509 100989
rect 156543 100961 156571 100989
rect 156357 92147 156385 92175
rect 156419 92147 156447 92175
rect 156481 92147 156509 92175
rect 156543 92147 156571 92175
rect 156357 92085 156385 92113
rect 156419 92085 156447 92113
rect 156481 92085 156509 92113
rect 156543 92085 156571 92113
rect 156357 92023 156385 92051
rect 156419 92023 156447 92051
rect 156481 92023 156509 92051
rect 156543 92023 156571 92051
rect 156357 91961 156385 91989
rect 156419 91961 156447 91989
rect 156481 91961 156509 91989
rect 156543 91961 156571 91989
rect 156357 83147 156385 83175
rect 156419 83147 156447 83175
rect 156481 83147 156509 83175
rect 156543 83147 156571 83175
rect 156357 83085 156385 83113
rect 156419 83085 156447 83113
rect 156481 83085 156509 83113
rect 156543 83085 156571 83113
rect 156357 83023 156385 83051
rect 156419 83023 156447 83051
rect 156481 83023 156509 83051
rect 156543 83023 156571 83051
rect 156357 82961 156385 82989
rect 156419 82961 156447 82989
rect 156481 82961 156509 82989
rect 156543 82961 156571 82989
rect 156357 74147 156385 74175
rect 156419 74147 156447 74175
rect 156481 74147 156509 74175
rect 156543 74147 156571 74175
rect 156357 74085 156385 74113
rect 156419 74085 156447 74113
rect 156481 74085 156509 74113
rect 156543 74085 156571 74113
rect 156357 74023 156385 74051
rect 156419 74023 156447 74051
rect 156481 74023 156509 74051
rect 156543 74023 156571 74051
rect 156357 73961 156385 73989
rect 156419 73961 156447 73989
rect 156481 73961 156509 73989
rect 156543 73961 156571 73989
rect 156357 65147 156385 65175
rect 156419 65147 156447 65175
rect 156481 65147 156509 65175
rect 156543 65147 156571 65175
rect 156357 65085 156385 65113
rect 156419 65085 156447 65113
rect 156481 65085 156509 65113
rect 156543 65085 156571 65113
rect 156357 65023 156385 65051
rect 156419 65023 156447 65051
rect 156481 65023 156509 65051
rect 156543 65023 156571 65051
rect 156357 64961 156385 64989
rect 156419 64961 156447 64989
rect 156481 64961 156509 64989
rect 156543 64961 156571 64989
rect 156357 56147 156385 56175
rect 156419 56147 156447 56175
rect 156481 56147 156509 56175
rect 156543 56147 156571 56175
rect 156357 56085 156385 56113
rect 156419 56085 156447 56113
rect 156481 56085 156509 56113
rect 156543 56085 156571 56113
rect 156357 56023 156385 56051
rect 156419 56023 156447 56051
rect 156481 56023 156509 56051
rect 156543 56023 156571 56051
rect 156357 55961 156385 55989
rect 156419 55961 156447 55989
rect 156481 55961 156509 55989
rect 156543 55961 156571 55989
rect 156357 47147 156385 47175
rect 156419 47147 156447 47175
rect 156481 47147 156509 47175
rect 156543 47147 156571 47175
rect 156357 47085 156385 47113
rect 156419 47085 156447 47113
rect 156481 47085 156509 47113
rect 156543 47085 156571 47113
rect 156357 47023 156385 47051
rect 156419 47023 156447 47051
rect 156481 47023 156509 47051
rect 156543 47023 156571 47051
rect 156357 46961 156385 46989
rect 156419 46961 156447 46989
rect 156481 46961 156509 46989
rect 156543 46961 156571 46989
rect 156357 38147 156385 38175
rect 156419 38147 156447 38175
rect 156481 38147 156509 38175
rect 156543 38147 156571 38175
rect 156357 38085 156385 38113
rect 156419 38085 156447 38113
rect 156481 38085 156509 38113
rect 156543 38085 156571 38113
rect 156357 38023 156385 38051
rect 156419 38023 156447 38051
rect 156481 38023 156509 38051
rect 156543 38023 156571 38051
rect 156357 37961 156385 37989
rect 156419 37961 156447 37989
rect 156481 37961 156509 37989
rect 156543 37961 156571 37989
rect 156357 29147 156385 29175
rect 156419 29147 156447 29175
rect 156481 29147 156509 29175
rect 156543 29147 156571 29175
rect 156357 29085 156385 29113
rect 156419 29085 156447 29113
rect 156481 29085 156509 29113
rect 156543 29085 156571 29113
rect 156357 29023 156385 29051
rect 156419 29023 156447 29051
rect 156481 29023 156509 29051
rect 156543 29023 156571 29051
rect 156357 28961 156385 28989
rect 156419 28961 156447 28989
rect 156481 28961 156509 28989
rect 156543 28961 156571 28989
rect 156357 20147 156385 20175
rect 156419 20147 156447 20175
rect 156481 20147 156509 20175
rect 156543 20147 156571 20175
rect 156357 20085 156385 20113
rect 156419 20085 156447 20113
rect 156481 20085 156509 20113
rect 156543 20085 156571 20113
rect 156357 20023 156385 20051
rect 156419 20023 156447 20051
rect 156481 20023 156509 20051
rect 156543 20023 156571 20051
rect 156357 19961 156385 19989
rect 156419 19961 156447 19989
rect 156481 19961 156509 19989
rect 156543 19961 156571 19989
rect 156357 11147 156385 11175
rect 156419 11147 156447 11175
rect 156481 11147 156509 11175
rect 156543 11147 156571 11175
rect 156357 11085 156385 11113
rect 156419 11085 156447 11113
rect 156481 11085 156509 11113
rect 156543 11085 156571 11113
rect 156357 11023 156385 11051
rect 156419 11023 156447 11051
rect 156481 11023 156509 11051
rect 156543 11023 156571 11051
rect 156357 10961 156385 10989
rect 156419 10961 156447 10989
rect 156481 10961 156509 10989
rect 156543 10961 156571 10989
rect 156357 2147 156385 2175
rect 156419 2147 156447 2175
rect 156481 2147 156509 2175
rect 156543 2147 156571 2175
rect 156357 2085 156385 2113
rect 156419 2085 156447 2113
rect 156481 2085 156509 2113
rect 156543 2085 156571 2113
rect 156357 2023 156385 2051
rect 156419 2023 156447 2051
rect 156481 2023 156509 2051
rect 156543 2023 156571 2051
rect 156357 1961 156385 1989
rect 156419 1961 156447 1989
rect 156481 1961 156509 1989
rect 156543 1961 156571 1989
rect 156357 -108 156385 -80
rect 156419 -108 156447 -80
rect 156481 -108 156509 -80
rect 156543 -108 156571 -80
rect 156357 -170 156385 -142
rect 156419 -170 156447 -142
rect 156481 -170 156509 -142
rect 156543 -170 156571 -142
rect 156357 -232 156385 -204
rect 156419 -232 156447 -204
rect 156481 -232 156509 -204
rect 156543 -232 156571 -204
rect 156357 -294 156385 -266
rect 156419 -294 156447 -266
rect 156481 -294 156509 -266
rect 156543 -294 156571 -266
rect 158217 130986 158245 131014
rect 158279 130986 158307 131014
rect 158341 130986 158369 131014
rect 158403 130986 158431 131014
rect 158217 130924 158245 130952
rect 158279 130924 158307 130952
rect 158341 130924 158369 130952
rect 158403 130924 158431 130952
rect 173577 130986 173605 131014
rect 173639 130986 173667 131014
rect 173701 130986 173729 131014
rect 173763 130986 173791 131014
rect 173577 130924 173605 130952
rect 173639 130924 173667 130952
rect 173701 130924 173729 130952
rect 173763 130924 173791 130952
rect 188937 130986 188965 131014
rect 188999 130986 189027 131014
rect 189061 130986 189089 131014
rect 189123 130986 189151 131014
rect 188937 130924 188965 130952
rect 188999 130924 189027 130952
rect 189061 130924 189089 130952
rect 189123 130924 189151 130952
rect 204297 131023 204325 131051
rect 204359 131023 204387 131051
rect 204421 131023 204449 131051
rect 204483 131023 204511 131051
rect 204297 130961 204325 130989
rect 204359 130961 204387 130989
rect 204421 130961 204449 130989
rect 204483 130961 204511 130989
rect 217797 128147 217825 128175
rect 217859 128147 217887 128175
rect 217921 128147 217949 128175
rect 217983 128147 218011 128175
rect 217797 128085 217825 128113
rect 217859 128085 217887 128113
rect 217921 128085 217949 128113
rect 217983 128085 218011 128113
rect 217797 128023 217825 128051
rect 217859 128023 217887 128051
rect 217921 128023 217949 128051
rect 217983 128023 218011 128051
rect 217797 127961 217825 127989
rect 217859 127961 217887 127989
rect 217921 127961 217949 127989
rect 217983 127961 218011 127989
rect 219657 299058 219685 299086
rect 219719 299058 219747 299086
rect 219781 299058 219809 299086
rect 219843 299058 219871 299086
rect 219657 298996 219685 299024
rect 219719 298996 219747 299024
rect 219781 298996 219809 299024
rect 219843 298996 219871 299024
rect 219657 298934 219685 298962
rect 219719 298934 219747 298962
rect 219781 298934 219809 298962
rect 219843 298934 219871 298962
rect 219657 298872 219685 298900
rect 219719 298872 219747 298900
rect 219781 298872 219809 298900
rect 219843 298872 219871 298900
rect 219657 293147 219685 293175
rect 219719 293147 219747 293175
rect 219781 293147 219809 293175
rect 219843 293147 219871 293175
rect 219657 293085 219685 293113
rect 219719 293085 219747 293113
rect 219781 293085 219809 293113
rect 219843 293085 219871 293113
rect 219657 293023 219685 293051
rect 219719 293023 219747 293051
rect 219781 293023 219809 293051
rect 219843 293023 219871 293051
rect 219657 292961 219685 292989
rect 219719 292961 219747 292989
rect 219781 292961 219809 292989
rect 219843 292961 219871 292989
rect 219657 284147 219685 284175
rect 219719 284147 219747 284175
rect 219781 284147 219809 284175
rect 219843 284147 219871 284175
rect 219657 284085 219685 284113
rect 219719 284085 219747 284113
rect 219781 284085 219809 284113
rect 219843 284085 219871 284113
rect 219657 284023 219685 284051
rect 219719 284023 219747 284051
rect 219781 284023 219809 284051
rect 219843 284023 219871 284051
rect 219657 283961 219685 283989
rect 219719 283961 219747 283989
rect 219781 283961 219809 283989
rect 219843 283961 219871 283989
rect 219657 275147 219685 275175
rect 219719 275147 219747 275175
rect 219781 275147 219809 275175
rect 219843 275147 219871 275175
rect 219657 275085 219685 275113
rect 219719 275085 219747 275113
rect 219781 275085 219809 275113
rect 219843 275085 219871 275113
rect 219657 275023 219685 275051
rect 219719 275023 219747 275051
rect 219781 275023 219809 275051
rect 219843 275023 219871 275051
rect 219657 274961 219685 274989
rect 219719 274961 219747 274989
rect 219781 274961 219809 274989
rect 219843 274961 219871 274989
rect 219657 266147 219685 266175
rect 219719 266147 219747 266175
rect 219781 266147 219809 266175
rect 219843 266147 219871 266175
rect 219657 266085 219685 266113
rect 219719 266085 219747 266113
rect 219781 266085 219809 266113
rect 219843 266085 219871 266113
rect 219657 266023 219685 266051
rect 219719 266023 219747 266051
rect 219781 266023 219809 266051
rect 219843 266023 219871 266051
rect 219657 265961 219685 265989
rect 219719 265961 219747 265989
rect 219781 265961 219809 265989
rect 219843 265961 219871 265989
rect 219657 257147 219685 257175
rect 219719 257147 219747 257175
rect 219781 257147 219809 257175
rect 219843 257147 219871 257175
rect 219657 257085 219685 257113
rect 219719 257085 219747 257113
rect 219781 257085 219809 257113
rect 219843 257085 219871 257113
rect 219657 257023 219685 257051
rect 219719 257023 219747 257051
rect 219781 257023 219809 257051
rect 219843 257023 219871 257051
rect 219657 256961 219685 256989
rect 219719 256961 219747 256989
rect 219781 256961 219809 256989
rect 219843 256961 219871 256989
rect 219657 248147 219685 248175
rect 219719 248147 219747 248175
rect 219781 248147 219809 248175
rect 219843 248147 219871 248175
rect 219657 248085 219685 248113
rect 219719 248085 219747 248113
rect 219781 248085 219809 248113
rect 219843 248085 219871 248113
rect 219657 248023 219685 248051
rect 219719 248023 219747 248051
rect 219781 248023 219809 248051
rect 219843 248023 219871 248051
rect 219657 247961 219685 247989
rect 219719 247961 219747 247989
rect 219781 247961 219809 247989
rect 219843 247961 219871 247989
rect 219657 239147 219685 239175
rect 219719 239147 219747 239175
rect 219781 239147 219809 239175
rect 219843 239147 219871 239175
rect 219657 239085 219685 239113
rect 219719 239085 219747 239113
rect 219781 239085 219809 239113
rect 219843 239085 219871 239113
rect 219657 239023 219685 239051
rect 219719 239023 219747 239051
rect 219781 239023 219809 239051
rect 219843 239023 219871 239051
rect 219657 238961 219685 238989
rect 219719 238961 219747 238989
rect 219781 238961 219809 238989
rect 219843 238961 219871 238989
rect 219657 230147 219685 230175
rect 219719 230147 219747 230175
rect 219781 230147 219809 230175
rect 219843 230147 219871 230175
rect 219657 230085 219685 230113
rect 219719 230085 219747 230113
rect 219781 230085 219809 230113
rect 219843 230085 219871 230113
rect 219657 230023 219685 230051
rect 219719 230023 219747 230051
rect 219781 230023 219809 230051
rect 219843 230023 219871 230051
rect 219657 229961 219685 229989
rect 219719 229961 219747 229989
rect 219781 229961 219809 229989
rect 219843 229961 219871 229989
rect 219657 221147 219685 221175
rect 219719 221147 219747 221175
rect 219781 221147 219809 221175
rect 219843 221147 219871 221175
rect 219657 221085 219685 221113
rect 219719 221085 219747 221113
rect 219781 221085 219809 221113
rect 219843 221085 219871 221113
rect 219657 221023 219685 221051
rect 219719 221023 219747 221051
rect 219781 221023 219809 221051
rect 219843 221023 219871 221051
rect 219657 220961 219685 220989
rect 219719 220961 219747 220989
rect 219781 220961 219809 220989
rect 219843 220961 219871 220989
rect 219657 212147 219685 212175
rect 219719 212147 219747 212175
rect 219781 212147 219809 212175
rect 219843 212147 219871 212175
rect 219657 212085 219685 212113
rect 219719 212085 219747 212113
rect 219781 212085 219809 212113
rect 219843 212085 219871 212113
rect 219657 212023 219685 212051
rect 219719 212023 219747 212051
rect 219781 212023 219809 212051
rect 219843 212023 219871 212051
rect 219657 211961 219685 211989
rect 219719 211961 219747 211989
rect 219781 211961 219809 211989
rect 219843 211961 219871 211989
rect 219657 203147 219685 203175
rect 219719 203147 219747 203175
rect 219781 203147 219809 203175
rect 219843 203147 219871 203175
rect 219657 203085 219685 203113
rect 219719 203085 219747 203113
rect 219781 203085 219809 203113
rect 219843 203085 219871 203113
rect 219657 203023 219685 203051
rect 219719 203023 219747 203051
rect 219781 203023 219809 203051
rect 219843 203023 219871 203051
rect 219657 202961 219685 202989
rect 219719 202961 219747 202989
rect 219781 202961 219809 202989
rect 219843 202961 219871 202989
rect 219657 194147 219685 194175
rect 219719 194147 219747 194175
rect 219781 194147 219809 194175
rect 219843 194147 219871 194175
rect 219657 194085 219685 194113
rect 219719 194085 219747 194113
rect 219781 194085 219809 194113
rect 219843 194085 219871 194113
rect 219657 194023 219685 194051
rect 219719 194023 219747 194051
rect 219781 194023 219809 194051
rect 219843 194023 219871 194051
rect 219657 193961 219685 193989
rect 219719 193961 219747 193989
rect 219781 193961 219809 193989
rect 219843 193961 219871 193989
rect 219657 185147 219685 185175
rect 219719 185147 219747 185175
rect 219781 185147 219809 185175
rect 219843 185147 219871 185175
rect 219657 185085 219685 185113
rect 219719 185085 219747 185113
rect 219781 185085 219809 185113
rect 219843 185085 219871 185113
rect 219657 185023 219685 185051
rect 219719 185023 219747 185051
rect 219781 185023 219809 185051
rect 219843 185023 219871 185051
rect 219657 184961 219685 184989
rect 219719 184961 219747 184989
rect 219781 184961 219809 184989
rect 219843 184961 219871 184989
rect 219657 176147 219685 176175
rect 219719 176147 219747 176175
rect 219781 176147 219809 176175
rect 219843 176147 219871 176175
rect 219657 176085 219685 176113
rect 219719 176085 219747 176113
rect 219781 176085 219809 176113
rect 219843 176085 219871 176113
rect 219657 176023 219685 176051
rect 219719 176023 219747 176051
rect 219781 176023 219809 176051
rect 219843 176023 219871 176051
rect 219657 175961 219685 175989
rect 219719 175961 219747 175989
rect 219781 175961 219809 175989
rect 219843 175961 219871 175989
rect 219657 167147 219685 167175
rect 219719 167147 219747 167175
rect 219781 167147 219809 167175
rect 219843 167147 219871 167175
rect 219657 167085 219685 167113
rect 219719 167085 219747 167113
rect 219781 167085 219809 167113
rect 219843 167085 219871 167113
rect 219657 167023 219685 167051
rect 219719 167023 219747 167051
rect 219781 167023 219809 167051
rect 219843 167023 219871 167051
rect 219657 166961 219685 166989
rect 219719 166961 219747 166989
rect 219781 166961 219809 166989
rect 219843 166961 219871 166989
rect 233157 298578 233185 298606
rect 233219 298578 233247 298606
rect 233281 298578 233309 298606
rect 233343 298578 233371 298606
rect 233157 298516 233185 298544
rect 233219 298516 233247 298544
rect 233281 298516 233309 298544
rect 233343 298516 233371 298544
rect 233157 298454 233185 298482
rect 233219 298454 233247 298482
rect 233281 298454 233309 298482
rect 233343 298454 233371 298482
rect 233157 298392 233185 298420
rect 233219 298392 233247 298420
rect 233281 298392 233309 298420
rect 233343 298392 233371 298420
rect 233157 290147 233185 290175
rect 233219 290147 233247 290175
rect 233281 290147 233309 290175
rect 233343 290147 233371 290175
rect 233157 290085 233185 290113
rect 233219 290085 233247 290113
rect 233281 290085 233309 290113
rect 233343 290085 233371 290113
rect 233157 290023 233185 290051
rect 233219 290023 233247 290051
rect 233281 290023 233309 290051
rect 233343 290023 233371 290051
rect 233157 289961 233185 289989
rect 233219 289961 233247 289989
rect 233281 289961 233309 289989
rect 233343 289961 233371 289989
rect 233157 281147 233185 281175
rect 233219 281147 233247 281175
rect 233281 281147 233309 281175
rect 233343 281147 233371 281175
rect 233157 281085 233185 281113
rect 233219 281085 233247 281113
rect 233281 281085 233309 281113
rect 233343 281085 233371 281113
rect 233157 281023 233185 281051
rect 233219 281023 233247 281051
rect 233281 281023 233309 281051
rect 233343 281023 233371 281051
rect 233157 280961 233185 280989
rect 233219 280961 233247 280989
rect 233281 280961 233309 280989
rect 233343 280961 233371 280989
rect 233157 272147 233185 272175
rect 233219 272147 233247 272175
rect 233281 272147 233309 272175
rect 233343 272147 233371 272175
rect 233157 272085 233185 272113
rect 233219 272085 233247 272113
rect 233281 272085 233309 272113
rect 233343 272085 233371 272113
rect 233157 272023 233185 272051
rect 233219 272023 233247 272051
rect 233281 272023 233309 272051
rect 233343 272023 233371 272051
rect 233157 271961 233185 271989
rect 233219 271961 233247 271989
rect 233281 271961 233309 271989
rect 233343 271961 233371 271989
rect 233157 263147 233185 263175
rect 233219 263147 233247 263175
rect 233281 263147 233309 263175
rect 233343 263147 233371 263175
rect 233157 263085 233185 263113
rect 233219 263085 233247 263113
rect 233281 263085 233309 263113
rect 233343 263085 233371 263113
rect 233157 263023 233185 263051
rect 233219 263023 233247 263051
rect 233281 263023 233309 263051
rect 233343 263023 233371 263051
rect 233157 262961 233185 262989
rect 233219 262961 233247 262989
rect 233281 262961 233309 262989
rect 233343 262961 233371 262989
rect 233157 254147 233185 254175
rect 233219 254147 233247 254175
rect 233281 254147 233309 254175
rect 233343 254147 233371 254175
rect 233157 254085 233185 254113
rect 233219 254085 233247 254113
rect 233281 254085 233309 254113
rect 233343 254085 233371 254113
rect 233157 254023 233185 254051
rect 233219 254023 233247 254051
rect 233281 254023 233309 254051
rect 233343 254023 233371 254051
rect 233157 253961 233185 253989
rect 233219 253961 233247 253989
rect 233281 253961 233309 253989
rect 233343 253961 233371 253989
rect 233157 245147 233185 245175
rect 233219 245147 233247 245175
rect 233281 245147 233309 245175
rect 233343 245147 233371 245175
rect 233157 245085 233185 245113
rect 233219 245085 233247 245113
rect 233281 245085 233309 245113
rect 233343 245085 233371 245113
rect 233157 245023 233185 245051
rect 233219 245023 233247 245051
rect 233281 245023 233309 245051
rect 233343 245023 233371 245051
rect 233157 244961 233185 244989
rect 233219 244961 233247 244989
rect 233281 244961 233309 244989
rect 233343 244961 233371 244989
rect 233157 236147 233185 236175
rect 233219 236147 233247 236175
rect 233281 236147 233309 236175
rect 233343 236147 233371 236175
rect 233157 236085 233185 236113
rect 233219 236085 233247 236113
rect 233281 236085 233309 236113
rect 233343 236085 233371 236113
rect 233157 236023 233185 236051
rect 233219 236023 233247 236051
rect 233281 236023 233309 236051
rect 233343 236023 233371 236051
rect 233157 235961 233185 235989
rect 233219 235961 233247 235989
rect 233281 235961 233309 235989
rect 233343 235961 233371 235989
rect 233157 227147 233185 227175
rect 233219 227147 233247 227175
rect 233281 227147 233309 227175
rect 233343 227147 233371 227175
rect 233157 227085 233185 227113
rect 233219 227085 233247 227113
rect 233281 227085 233309 227113
rect 233343 227085 233371 227113
rect 233157 227023 233185 227051
rect 233219 227023 233247 227051
rect 233281 227023 233309 227051
rect 233343 227023 233371 227051
rect 233157 226961 233185 226989
rect 233219 226961 233247 226989
rect 233281 226961 233309 226989
rect 233343 226961 233371 226989
rect 233157 218147 233185 218175
rect 233219 218147 233247 218175
rect 233281 218147 233309 218175
rect 233343 218147 233371 218175
rect 233157 218085 233185 218113
rect 233219 218085 233247 218113
rect 233281 218085 233309 218113
rect 233343 218085 233371 218113
rect 233157 218023 233185 218051
rect 233219 218023 233247 218051
rect 233281 218023 233309 218051
rect 233343 218023 233371 218051
rect 233157 217961 233185 217989
rect 233219 217961 233247 217989
rect 233281 217961 233309 217989
rect 233343 217961 233371 217989
rect 233157 209147 233185 209175
rect 233219 209147 233247 209175
rect 233281 209147 233309 209175
rect 233343 209147 233371 209175
rect 233157 209085 233185 209113
rect 233219 209085 233247 209113
rect 233281 209085 233309 209113
rect 233343 209085 233371 209113
rect 233157 209023 233185 209051
rect 233219 209023 233247 209051
rect 233281 209023 233309 209051
rect 233343 209023 233371 209051
rect 233157 208961 233185 208989
rect 233219 208961 233247 208989
rect 233281 208961 233309 208989
rect 233343 208961 233371 208989
rect 233157 200147 233185 200175
rect 233219 200147 233247 200175
rect 233281 200147 233309 200175
rect 233343 200147 233371 200175
rect 233157 200085 233185 200113
rect 233219 200085 233247 200113
rect 233281 200085 233309 200113
rect 233343 200085 233371 200113
rect 233157 200023 233185 200051
rect 233219 200023 233247 200051
rect 233281 200023 233309 200051
rect 233343 200023 233371 200051
rect 233157 199961 233185 199989
rect 233219 199961 233247 199989
rect 233281 199961 233309 199989
rect 233343 199961 233371 199989
rect 233157 191147 233185 191175
rect 233219 191147 233247 191175
rect 233281 191147 233309 191175
rect 233343 191147 233371 191175
rect 233157 191085 233185 191113
rect 233219 191085 233247 191113
rect 233281 191085 233309 191113
rect 233343 191085 233371 191113
rect 233157 191023 233185 191051
rect 233219 191023 233247 191051
rect 233281 191023 233309 191051
rect 233343 191023 233371 191051
rect 233157 190961 233185 190989
rect 233219 190961 233247 190989
rect 233281 190961 233309 190989
rect 233343 190961 233371 190989
rect 233157 182147 233185 182175
rect 233219 182147 233247 182175
rect 233281 182147 233309 182175
rect 233343 182147 233371 182175
rect 233157 182085 233185 182113
rect 233219 182085 233247 182113
rect 233281 182085 233309 182113
rect 233343 182085 233371 182113
rect 233157 182023 233185 182051
rect 233219 182023 233247 182051
rect 233281 182023 233309 182051
rect 233343 182023 233371 182051
rect 233157 181961 233185 181989
rect 233219 181961 233247 181989
rect 233281 181961 233309 181989
rect 233343 181961 233371 181989
rect 233157 173147 233185 173175
rect 233219 173147 233247 173175
rect 233281 173147 233309 173175
rect 233343 173147 233371 173175
rect 233157 173085 233185 173113
rect 233219 173085 233247 173113
rect 233281 173085 233309 173113
rect 233343 173085 233371 173113
rect 233157 173023 233185 173051
rect 233219 173023 233247 173051
rect 233281 173023 233309 173051
rect 233343 173023 233371 173051
rect 233157 172961 233185 172989
rect 233219 172961 233247 172989
rect 233281 172961 233309 172989
rect 233343 172961 233371 172989
rect 233157 164147 233185 164175
rect 233219 164147 233247 164175
rect 233281 164147 233309 164175
rect 233343 164147 233371 164175
rect 233157 164085 233185 164113
rect 233219 164085 233247 164113
rect 233281 164085 233309 164113
rect 233343 164085 233371 164113
rect 233157 164023 233185 164051
rect 233219 164023 233247 164051
rect 233281 164023 233309 164051
rect 233343 164023 233371 164051
rect 233157 163961 233185 163989
rect 233219 163961 233247 163989
rect 233281 163961 233309 163989
rect 233343 163961 233371 163989
rect 219657 158147 219685 158175
rect 219719 158147 219747 158175
rect 219781 158147 219809 158175
rect 219843 158147 219871 158175
rect 219657 158085 219685 158113
rect 219719 158085 219747 158113
rect 219781 158085 219809 158113
rect 219843 158085 219871 158113
rect 219657 158023 219685 158051
rect 219719 158023 219747 158051
rect 219781 158023 219809 158051
rect 219843 158023 219871 158051
rect 219657 157961 219685 157989
rect 219719 157961 219747 157989
rect 219781 157961 219809 157989
rect 219843 157961 219871 157989
rect 224259 158147 224287 158175
rect 224321 158147 224349 158175
rect 224259 158085 224287 158113
rect 224321 158085 224349 158113
rect 224259 158023 224287 158051
rect 224321 158023 224349 158051
rect 224259 157961 224287 157989
rect 224321 157961 224349 157989
rect 231939 155147 231967 155175
rect 232001 155147 232029 155175
rect 231939 155085 231967 155113
rect 232001 155085 232029 155113
rect 231939 155023 231967 155051
rect 232001 155023 232029 155051
rect 231939 154961 231967 154989
rect 232001 154961 232029 154989
rect 233157 155147 233185 155175
rect 233219 155147 233247 155175
rect 233281 155147 233309 155175
rect 233343 155147 233371 155175
rect 233157 155085 233185 155113
rect 233219 155085 233247 155113
rect 233281 155085 233309 155113
rect 233343 155085 233371 155113
rect 233157 155023 233185 155051
rect 233219 155023 233247 155051
rect 233281 155023 233309 155051
rect 233343 155023 233371 155051
rect 233157 154961 233185 154989
rect 233219 154961 233247 154989
rect 233281 154961 233309 154989
rect 233343 154961 233371 154989
rect 219657 149147 219685 149175
rect 219719 149147 219747 149175
rect 219781 149147 219809 149175
rect 219843 149147 219871 149175
rect 219657 149085 219685 149113
rect 219719 149085 219747 149113
rect 219781 149085 219809 149113
rect 219843 149085 219871 149113
rect 219657 149023 219685 149051
rect 219719 149023 219747 149051
rect 219781 149023 219809 149051
rect 219843 149023 219871 149051
rect 219657 148961 219685 148989
rect 219719 148961 219747 148989
rect 219781 148961 219809 148989
rect 219843 148961 219871 148989
rect 224259 149147 224287 149175
rect 224321 149147 224349 149175
rect 224259 149085 224287 149113
rect 224321 149085 224349 149113
rect 224259 149023 224287 149051
rect 224321 149023 224349 149051
rect 224259 148961 224287 148989
rect 224321 148961 224349 148989
rect 231939 146147 231967 146175
rect 232001 146147 232029 146175
rect 231939 146085 231967 146113
rect 232001 146085 232029 146113
rect 231939 146023 231967 146051
rect 232001 146023 232029 146051
rect 231939 145961 231967 145989
rect 232001 145961 232029 145989
rect 233157 146147 233185 146175
rect 233219 146147 233247 146175
rect 233281 146147 233309 146175
rect 233343 146147 233371 146175
rect 233157 146085 233185 146113
rect 233219 146085 233247 146113
rect 233281 146085 233309 146113
rect 233343 146085 233371 146113
rect 233157 146023 233185 146051
rect 233219 146023 233247 146051
rect 233281 146023 233309 146051
rect 233343 146023 233371 146051
rect 233157 145961 233185 145989
rect 233219 145961 233247 145989
rect 233281 145961 233309 145989
rect 233343 145961 233371 145989
rect 219657 140147 219685 140175
rect 219719 140147 219747 140175
rect 219781 140147 219809 140175
rect 219843 140147 219871 140175
rect 219657 140085 219685 140113
rect 219719 140085 219747 140113
rect 219781 140085 219809 140113
rect 219843 140085 219871 140113
rect 219657 140023 219685 140051
rect 219719 140023 219747 140051
rect 219781 140023 219809 140051
rect 219843 140023 219871 140051
rect 219657 139961 219685 139989
rect 219719 139961 219747 139989
rect 219781 139961 219809 139989
rect 219843 139961 219871 139989
rect 224259 140147 224287 140175
rect 224321 140147 224349 140175
rect 224259 140085 224287 140113
rect 224321 140085 224349 140113
rect 224259 140023 224287 140051
rect 224321 140023 224349 140051
rect 224259 139961 224287 139989
rect 224321 139961 224349 139989
rect 231939 137147 231967 137175
rect 232001 137147 232029 137175
rect 231939 137085 231967 137113
rect 232001 137085 232029 137113
rect 231939 137023 231967 137051
rect 232001 137023 232029 137051
rect 231939 136961 231967 136989
rect 232001 136961 232029 136989
rect 233157 137147 233185 137175
rect 233219 137147 233247 137175
rect 233281 137147 233309 137175
rect 233343 137147 233371 137175
rect 233157 137085 233185 137113
rect 233219 137085 233247 137113
rect 233281 137085 233309 137113
rect 233343 137085 233371 137113
rect 233157 137023 233185 137051
rect 233219 137023 233247 137051
rect 233281 137023 233309 137051
rect 233343 137023 233371 137051
rect 233157 136961 233185 136989
rect 233219 136961 233247 136989
rect 233281 136961 233309 136989
rect 233343 136961 233371 136989
rect 219657 131147 219685 131175
rect 219719 131147 219747 131175
rect 219781 131147 219809 131175
rect 219843 131147 219871 131175
rect 219657 131085 219685 131113
rect 219719 131085 219747 131113
rect 219781 131085 219809 131113
rect 219843 131085 219871 131113
rect 219657 131023 219685 131051
rect 219719 131023 219747 131051
rect 219781 131023 219809 131051
rect 219843 131023 219871 131051
rect 219657 130961 219685 130989
rect 219719 130961 219747 130989
rect 219781 130961 219809 130989
rect 219843 130961 219871 130989
rect 233157 128147 233185 128175
rect 233219 128147 233247 128175
rect 233281 128147 233309 128175
rect 233343 128147 233371 128175
rect 233157 128085 233185 128113
rect 233219 128085 233247 128113
rect 233281 128085 233309 128113
rect 233343 128085 233371 128113
rect 233157 128023 233185 128051
rect 233219 128023 233247 128051
rect 233281 128023 233309 128051
rect 233343 128023 233371 128051
rect 233157 127961 233185 127989
rect 233219 127961 233247 127989
rect 233281 127961 233309 127989
rect 233343 127961 233371 127989
rect 235017 299058 235045 299086
rect 235079 299058 235107 299086
rect 235141 299058 235169 299086
rect 235203 299058 235231 299086
rect 235017 298996 235045 299024
rect 235079 298996 235107 299024
rect 235141 298996 235169 299024
rect 235203 298996 235231 299024
rect 235017 298934 235045 298962
rect 235079 298934 235107 298962
rect 235141 298934 235169 298962
rect 235203 298934 235231 298962
rect 235017 298872 235045 298900
rect 235079 298872 235107 298900
rect 235141 298872 235169 298900
rect 235203 298872 235231 298900
rect 235017 293147 235045 293175
rect 235079 293147 235107 293175
rect 235141 293147 235169 293175
rect 235203 293147 235231 293175
rect 235017 293085 235045 293113
rect 235079 293085 235107 293113
rect 235141 293085 235169 293113
rect 235203 293085 235231 293113
rect 235017 293023 235045 293051
rect 235079 293023 235107 293051
rect 235141 293023 235169 293051
rect 235203 293023 235231 293051
rect 235017 292961 235045 292989
rect 235079 292961 235107 292989
rect 235141 292961 235169 292989
rect 235203 292961 235231 292989
rect 235017 284147 235045 284175
rect 235079 284147 235107 284175
rect 235141 284147 235169 284175
rect 235203 284147 235231 284175
rect 235017 284085 235045 284113
rect 235079 284085 235107 284113
rect 235141 284085 235169 284113
rect 235203 284085 235231 284113
rect 235017 284023 235045 284051
rect 235079 284023 235107 284051
rect 235141 284023 235169 284051
rect 235203 284023 235231 284051
rect 235017 283961 235045 283989
rect 235079 283961 235107 283989
rect 235141 283961 235169 283989
rect 235203 283961 235231 283989
rect 235017 275147 235045 275175
rect 235079 275147 235107 275175
rect 235141 275147 235169 275175
rect 235203 275147 235231 275175
rect 235017 275085 235045 275113
rect 235079 275085 235107 275113
rect 235141 275085 235169 275113
rect 235203 275085 235231 275113
rect 235017 275023 235045 275051
rect 235079 275023 235107 275051
rect 235141 275023 235169 275051
rect 235203 275023 235231 275051
rect 235017 274961 235045 274989
rect 235079 274961 235107 274989
rect 235141 274961 235169 274989
rect 235203 274961 235231 274989
rect 235017 266147 235045 266175
rect 235079 266147 235107 266175
rect 235141 266147 235169 266175
rect 235203 266147 235231 266175
rect 235017 266085 235045 266113
rect 235079 266085 235107 266113
rect 235141 266085 235169 266113
rect 235203 266085 235231 266113
rect 235017 266023 235045 266051
rect 235079 266023 235107 266051
rect 235141 266023 235169 266051
rect 235203 266023 235231 266051
rect 235017 265961 235045 265989
rect 235079 265961 235107 265989
rect 235141 265961 235169 265989
rect 235203 265961 235231 265989
rect 235017 257147 235045 257175
rect 235079 257147 235107 257175
rect 235141 257147 235169 257175
rect 235203 257147 235231 257175
rect 235017 257085 235045 257113
rect 235079 257085 235107 257113
rect 235141 257085 235169 257113
rect 235203 257085 235231 257113
rect 235017 257023 235045 257051
rect 235079 257023 235107 257051
rect 235141 257023 235169 257051
rect 235203 257023 235231 257051
rect 235017 256961 235045 256989
rect 235079 256961 235107 256989
rect 235141 256961 235169 256989
rect 235203 256961 235231 256989
rect 235017 248147 235045 248175
rect 235079 248147 235107 248175
rect 235141 248147 235169 248175
rect 235203 248147 235231 248175
rect 235017 248085 235045 248113
rect 235079 248085 235107 248113
rect 235141 248085 235169 248113
rect 235203 248085 235231 248113
rect 235017 248023 235045 248051
rect 235079 248023 235107 248051
rect 235141 248023 235169 248051
rect 235203 248023 235231 248051
rect 235017 247961 235045 247989
rect 235079 247961 235107 247989
rect 235141 247961 235169 247989
rect 235203 247961 235231 247989
rect 235017 239147 235045 239175
rect 235079 239147 235107 239175
rect 235141 239147 235169 239175
rect 235203 239147 235231 239175
rect 235017 239085 235045 239113
rect 235079 239085 235107 239113
rect 235141 239085 235169 239113
rect 235203 239085 235231 239113
rect 235017 239023 235045 239051
rect 235079 239023 235107 239051
rect 235141 239023 235169 239051
rect 235203 239023 235231 239051
rect 235017 238961 235045 238989
rect 235079 238961 235107 238989
rect 235141 238961 235169 238989
rect 235203 238961 235231 238989
rect 235017 230147 235045 230175
rect 235079 230147 235107 230175
rect 235141 230147 235169 230175
rect 235203 230147 235231 230175
rect 235017 230085 235045 230113
rect 235079 230085 235107 230113
rect 235141 230085 235169 230113
rect 235203 230085 235231 230113
rect 235017 230023 235045 230051
rect 235079 230023 235107 230051
rect 235141 230023 235169 230051
rect 235203 230023 235231 230051
rect 235017 229961 235045 229989
rect 235079 229961 235107 229989
rect 235141 229961 235169 229989
rect 235203 229961 235231 229989
rect 235017 221147 235045 221175
rect 235079 221147 235107 221175
rect 235141 221147 235169 221175
rect 235203 221147 235231 221175
rect 235017 221085 235045 221113
rect 235079 221085 235107 221113
rect 235141 221085 235169 221113
rect 235203 221085 235231 221113
rect 235017 221023 235045 221051
rect 235079 221023 235107 221051
rect 235141 221023 235169 221051
rect 235203 221023 235231 221051
rect 235017 220961 235045 220989
rect 235079 220961 235107 220989
rect 235141 220961 235169 220989
rect 235203 220961 235231 220989
rect 235017 212147 235045 212175
rect 235079 212147 235107 212175
rect 235141 212147 235169 212175
rect 235203 212147 235231 212175
rect 235017 212085 235045 212113
rect 235079 212085 235107 212113
rect 235141 212085 235169 212113
rect 235203 212085 235231 212113
rect 235017 212023 235045 212051
rect 235079 212023 235107 212051
rect 235141 212023 235169 212051
rect 235203 212023 235231 212051
rect 235017 211961 235045 211989
rect 235079 211961 235107 211989
rect 235141 211961 235169 211989
rect 235203 211961 235231 211989
rect 235017 203147 235045 203175
rect 235079 203147 235107 203175
rect 235141 203147 235169 203175
rect 235203 203147 235231 203175
rect 235017 203085 235045 203113
rect 235079 203085 235107 203113
rect 235141 203085 235169 203113
rect 235203 203085 235231 203113
rect 235017 203023 235045 203051
rect 235079 203023 235107 203051
rect 235141 203023 235169 203051
rect 235203 203023 235231 203051
rect 235017 202961 235045 202989
rect 235079 202961 235107 202989
rect 235141 202961 235169 202989
rect 235203 202961 235231 202989
rect 235017 194147 235045 194175
rect 235079 194147 235107 194175
rect 235141 194147 235169 194175
rect 235203 194147 235231 194175
rect 235017 194085 235045 194113
rect 235079 194085 235107 194113
rect 235141 194085 235169 194113
rect 235203 194085 235231 194113
rect 235017 194023 235045 194051
rect 235079 194023 235107 194051
rect 235141 194023 235169 194051
rect 235203 194023 235231 194051
rect 235017 193961 235045 193989
rect 235079 193961 235107 193989
rect 235141 193961 235169 193989
rect 235203 193961 235231 193989
rect 248517 298578 248545 298606
rect 248579 298578 248607 298606
rect 248641 298578 248669 298606
rect 248703 298578 248731 298606
rect 248517 298516 248545 298544
rect 248579 298516 248607 298544
rect 248641 298516 248669 298544
rect 248703 298516 248731 298544
rect 248517 298454 248545 298482
rect 248579 298454 248607 298482
rect 248641 298454 248669 298482
rect 248703 298454 248731 298482
rect 248517 298392 248545 298420
rect 248579 298392 248607 298420
rect 248641 298392 248669 298420
rect 248703 298392 248731 298420
rect 248517 290147 248545 290175
rect 248579 290147 248607 290175
rect 248641 290147 248669 290175
rect 248703 290147 248731 290175
rect 248517 290085 248545 290113
rect 248579 290085 248607 290113
rect 248641 290085 248669 290113
rect 248703 290085 248731 290113
rect 248517 290023 248545 290051
rect 248579 290023 248607 290051
rect 248641 290023 248669 290051
rect 248703 290023 248731 290051
rect 248517 289961 248545 289989
rect 248579 289961 248607 289989
rect 248641 289961 248669 289989
rect 248703 289961 248731 289989
rect 248517 281147 248545 281175
rect 248579 281147 248607 281175
rect 248641 281147 248669 281175
rect 248703 281147 248731 281175
rect 248517 281085 248545 281113
rect 248579 281085 248607 281113
rect 248641 281085 248669 281113
rect 248703 281085 248731 281113
rect 248517 281023 248545 281051
rect 248579 281023 248607 281051
rect 248641 281023 248669 281051
rect 248703 281023 248731 281051
rect 248517 280961 248545 280989
rect 248579 280961 248607 280989
rect 248641 280961 248669 280989
rect 248703 280961 248731 280989
rect 248517 272147 248545 272175
rect 248579 272147 248607 272175
rect 248641 272147 248669 272175
rect 248703 272147 248731 272175
rect 248517 272085 248545 272113
rect 248579 272085 248607 272113
rect 248641 272085 248669 272113
rect 248703 272085 248731 272113
rect 248517 272023 248545 272051
rect 248579 272023 248607 272051
rect 248641 272023 248669 272051
rect 248703 272023 248731 272051
rect 248517 271961 248545 271989
rect 248579 271961 248607 271989
rect 248641 271961 248669 271989
rect 248703 271961 248731 271989
rect 248517 263147 248545 263175
rect 248579 263147 248607 263175
rect 248641 263147 248669 263175
rect 248703 263147 248731 263175
rect 248517 263085 248545 263113
rect 248579 263085 248607 263113
rect 248641 263085 248669 263113
rect 248703 263085 248731 263113
rect 248517 263023 248545 263051
rect 248579 263023 248607 263051
rect 248641 263023 248669 263051
rect 248703 263023 248731 263051
rect 248517 262961 248545 262989
rect 248579 262961 248607 262989
rect 248641 262961 248669 262989
rect 248703 262961 248731 262989
rect 248517 254147 248545 254175
rect 248579 254147 248607 254175
rect 248641 254147 248669 254175
rect 248703 254147 248731 254175
rect 248517 254085 248545 254113
rect 248579 254085 248607 254113
rect 248641 254085 248669 254113
rect 248703 254085 248731 254113
rect 248517 254023 248545 254051
rect 248579 254023 248607 254051
rect 248641 254023 248669 254051
rect 248703 254023 248731 254051
rect 248517 253961 248545 253989
rect 248579 253961 248607 253989
rect 248641 253961 248669 253989
rect 248703 253961 248731 253989
rect 248517 245147 248545 245175
rect 248579 245147 248607 245175
rect 248641 245147 248669 245175
rect 248703 245147 248731 245175
rect 248517 245085 248545 245113
rect 248579 245085 248607 245113
rect 248641 245085 248669 245113
rect 248703 245085 248731 245113
rect 248517 245023 248545 245051
rect 248579 245023 248607 245051
rect 248641 245023 248669 245051
rect 248703 245023 248731 245051
rect 248517 244961 248545 244989
rect 248579 244961 248607 244989
rect 248641 244961 248669 244989
rect 248703 244961 248731 244989
rect 248517 236147 248545 236175
rect 248579 236147 248607 236175
rect 248641 236147 248669 236175
rect 248703 236147 248731 236175
rect 248517 236085 248545 236113
rect 248579 236085 248607 236113
rect 248641 236085 248669 236113
rect 248703 236085 248731 236113
rect 248517 236023 248545 236051
rect 248579 236023 248607 236051
rect 248641 236023 248669 236051
rect 248703 236023 248731 236051
rect 248517 235961 248545 235989
rect 248579 235961 248607 235989
rect 248641 235961 248669 235989
rect 248703 235961 248731 235989
rect 248517 227147 248545 227175
rect 248579 227147 248607 227175
rect 248641 227147 248669 227175
rect 248703 227147 248731 227175
rect 248517 227085 248545 227113
rect 248579 227085 248607 227113
rect 248641 227085 248669 227113
rect 248703 227085 248731 227113
rect 248517 227023 248545 227051
rect 248579 227023 248607 227051
rect 248641 227023 248669 227051
rect 248703 227023 248731 227051
rect 248517 226961 248545 226989
rect 248579 226961 248607 226989
rect 248641 226961 248669 226989
rect 248703 226961 248731 226989
rect 248517 218147 248545 218175
rect 248579 218147 248607 218175
rect 248641 218147 248669 218175
rect 248703 218147 248731 218175
rect 248517 218085 248545 218113
rect 248579 218085 248607 218113
rect 248641 218085 248669 218113
rect 248703 218085 248731 218113
rect 248517 218023 248545 218051
rect 248579 218023 248607 218051
rect 248641 218023 248669 218051
rect 248703 218023 248731 218051
rect 248517 217961 248545 217989
rect 248579 217961 248607 217989
rect 248641 217961 248669 217989
rect 248703 217961 248731 217989
rect 248517 209147 248545 209175
rect 248579 209147 248607 209175
rect 248641 209147 248669 209175
rect 248703 209147 248731 209175
rect 248517 209085 248545 209113
rect 248579 209085 248607 209113
rect 248641 209085 248669 209113
rect 248703 209085 248731 209113
rect 248517 209023 248545 209051
rect 248579 209023 248607 209051
rect 248641 209023 248669 209051
rect 248703 209023 248731 209051
rect 248517 208961 248545 208989
rect 248579 208961 248607 208989
rect 248641 208961 248669 208989
rect 248703 208961 248731 208989
rect 248517 200147 248545 200175
rect 248579 200147 248607 200175
rect 248641 200147 248669 200175
rect 248703 200147 248731 200175
rect 248517 200085 248545 200113
rect 248579 200085 248607 200113
rect 248641 200085 248669 200113
rect 248703 200085 248731 200113
rect 248517 200023 248545 200051
rect 248579 200023 248607 200051
rect 248641 200023 248669 200051
rect 248703 200023 248731 200051
rect 248517 199961 248545 199989
rect 248579 199961 248607 199989
rect 248641 199961 248669 199989
rect 248703 199961 248731 199989
rect 248517 191147 248545 191175
rect 248579 191147 248607 191175
rect 248641 191147 248669 191175
rect 248703 191147 248731 191175
rect 248517 191085 248545 191113
rect 248579 191085 248607 191113
rect 248641 191085 248669 191113
rect 248703 191085 248731 191113
rect 248517 191023 248545 191051
rect 248579 191023 248607 191051
rect 248641 191023 248669 191051
rect 248703 191023 248731 191051
rect 248517 190961 248545 190989
rect 248579 190961 248607 190989
rect 248641 190961 248669 190989
rect 248703 190961 248731 190989
rect 250377 299058 250405 299086
rect 250439 299058 250467 299086
rect 250501 299058 250529 299086
rect 250563 299058 250591 299086
rect 250377 298996 250405 299024
rect 250439 298996 250467 299024
rect 250501 298996 250529 299024
rect 250563 298996 250591 299024
rect 250377 298934 250405 298962
rect 250439 298934 250467 298962
rect 250501 298934 250529 298962
rect 250563 298934 250591 298962
rect 250377 298872 250405 298900
rect 250439 298872 250467 298900
rect 250501 298872 250529 298900
rect 250563 298872 250591 298900
rect 250377 293147 250405 293175
rect 250439 293147 250467 293175
rect 250501 293147 250529 293175
rect 250563 293147 250591 293175
rect 250377 293085 250405 293113
rect 250439 293085 250467 293113
rect 250501 293085 250529 293113
rect 250563 293085 250591 293113
rect 250377 293023 250405 293051
rect 250439 293023 250467 293051
rect 250501 293023 250529 293051
rect 250563 293023 250591 293051
rect 250377 292961 250405 292989
rect 250439 292961 250467 292989
rect 250501 292961 250529 292989
rect 250563 292961 250591 292989
rect 250377 284147 250405 284175
rect 250439 284147 250467 284175
rect 250501 284147 250529 284175
rect 250563 284147 250591 284175
rect 250377 284085 250405 284113
rect 250439 284085 250467 284113
rect 250501 284085 250529 284113
rect 250563 284085 250591 284113
rect 250377 284023 250405 284051
rect 250439 284023 250467 284051
rect 250501 284023 250529 284051
rect 250563 284023 250591 284051
rect 250377 283961 250405 283989
rect 250439 283961 250467 283989
rect 250501 283961 250529 283989
rect 250563 283961 250591 283989
rect 250377 275147 250405 275175
rect 250439 275147 250467 275175
rect 250501 275147 250529 275175
rect 250563 275147 250591 275175
rect 250377 275085 250405 275113
rect 250439 275085 250467 275113
rect 250501 275085 250529 275113
rect 250563 275085 250591 275113
rect 250377 275023 250405 275051
rect 250439 275023 250467 275051
rect 250501 275023 250529 275051
rect 250563 275023 250591 275051
rect 250377 274961 250405 274989
rect 250439 274961 250467 274989
rect 250501 274961 250529 274989
rect 250563 274961 250591 274989
rect 250377 266147 250405 266175
rect 250439 266147 250467 266175
rect 250501 266147 250529 266175
rect 250563 266147 250591 266175
rect 250377 266085 250405 266113
rect 250439 266085 250467 266113
rect 250501 266085 250529 266113
rect 250563 266085 250591 266113
rect 250377 266023 250405 266051
rect 250439 266023 250467 266051
rect 250501 266023 250529 266051
rect 250563 266023 250591 266051
rect 250377 265961 250405 265989
rect 250439 265961 250467 265989
rect 250501 265961 250529 265989
rect 250563 265961 250591 265989
rect 250377 257147 250405 257175
rect 250439 257147 250467 257175
rect 250501 257147 250529 257175
rect 250563 257147 250591 257175
rect 250377 257085 250405 257113
rect 250439 257085 250467 257113
rect 250501 257085 250529 257113
rect 250563 257085 250591 257113
rect 250377 257023 250405 257051
rect 250439 257023 250467 257051
rect 250501 257023 250529 257051
rect 250563 257023 250591 257051
rect 250377 256961 250405 256989
rect 250439 256961 250467 256989
rect 250501 256961 250529 256989
rect 250563 256961 250591 256989
rect 250377 248147 250405 248175
rect 250439 248147 250467 248175
rect 250501 248147 250529 248175
rect 250563 248147 250591 248175
rect 250377 248085 250405 248113
rect 250439 248085 250467 248113
rect 250501 248085 250529 248113
rect 250563 248085 250591 248113
rect 250377 248023 250405 248051
rect 250439 248023 250467 248051
rect 250501 248023 250529 248051
rect 250563 248023 250591 248051
rect 250377 247961 250405 247989
rect 250439 247961 250467 247989
rect 250501 247961 250529 247989
rect 250563 247961 250591 247989
rect 250377 239147 250405 239175
rect 250439 239147 250467 239175
rect 250501 239147 250529 239175
rect 250563 239147 250591 239175
rect 250377 239085 250405 239113
rect 250439 239085 250467 239113
rect 250501 239085 250529 239113
rect 250563 239085 250591 239113
rect 250377 239023 250405 239051
rect 250439 239023 250467 239051
rect 250501 239023 250529 239051
rect 250563 239023 250591 239051
rect 250377 238961 250405 238989
rect 250439 238961 250467 238989
rect 250501 238961 250529 238989
rect 250563 238961 250591 238989
rect 250377 230147 250405 230175
rect 250439 230147 250467 230175
rect 250501 230147 250529 230175
rect 250563 230147 250591 230175
rect 250377 230085 250405 230113
rect 250439 230085 250467 230113
rect 250501 230085 250529 230113
rect 250563 230085 250591 230113
rect 250377 230023 250405 230051
rect 250439 230023 250467 230051
rect 250501 230023 250529 230051
rect 250563 230023 250591 230051
rect 250377 229961 250405 229989
rect 250439 229961 250467 229989
rect 250501 229961 250529 229989
rect 250563 229961 250591 229989
rect 250377 221147 250405 221175
rect 250439 221147 250467 221175
rect 250501 221147 250529 221175
rect 250563 221147 250591 221175
rect 250377 221085 250405 221113
rect 250439 221085 250467 221113
rect 250501 221085 250529 221113
rect 250563 221085 250591 221113
rect 250377 221023 250405 221051
rect 250439 221023 250467 221051
rect 250501 221023 250529 221051
rect 250563 221023 250591 221051
rect 250377 220961 250405 220989
rect 250439 220961 250467 220989
rect 250501 220961 250529 220989
rect 250563 220961 250591 220989
rect 250377 212147 250405 212175
rect 250439 212147 250467 212175
rect 250501 212147 250529 212175
rect 250563 212147 250591 212175
rect 250377 212085 250405 212113
rect 250439 212085 250467 212113
rect 250501 212085 250529 212113
rect 250563 212085 250591 212113
rect 250377 212023 250405 212051
rect 250439 212023 250467 212051
rect 250501 212023 250529 212051
rect 250563 212023 250591 212051
rect 250377 211961 250405 211989
rect 250439 211961 250467 211989
rect 250501 211961 250529 211989
rect 250563 211961 250591 211989
rect 250377 203147 250405 203175
rect 250439 203147 250467 203175
rect 250501 203147 250529 203175
rect 250563 203147 250591 203175
rect 250377 203085 250405 203113
rect 250439 203085 250467 203113
rect 250501 203085 250529 203113
rect 250563 203085 250591 203113
rect 250377 203023 250405 203051
rect 250439 203023 250467 203051
rect 250501 203023 250529 203051
rect 250563 203023 250591 203051
rect 250377 202961 250405 202989
rect 250439 202961 250467 202989
rect 250501 202961 250529 202989
rect 250563 202961 250591 202989
rect 250377 194147 250405 194175
rect 250439 194147 250467 194175
rect 250501 194147 250529 194175
rect 250563 194147 250591 194175
rect 250377 194085 250405 194113
rect 250439 194085 250467 194113
rect 250501 194085 250529 194113
rect 250563 194085 250591 194113
rect 250377 194023 250405 194051
rect 250439 194023 250467 194051
rect 250501 194023 250529 194051
rect 250563 194023 250591 194051
rect 250377 193961 250405 193989
rect 250439 193961 250467 193989
rect 250501 193961 250529 193989
rect 250563 193961 250591 193989
rect 263877 298578 263905 298606
rect 263939 298578 263967 298606
rect 264001 298578 264029 298606
rect 264063 298578 264091 298606
rect 263877 298516 263905 298544
rect 263939 298516 263967 298544
rect 264001 298516 264029 298544
rect 264063 298516 264091 298544
rect 263877 298454 263905 298482
rect 263939 298454 263967 298482
rect 264001 298454 264029 298482
rect 264063 298454 264091 298482
rect 263877 298392 263905 298420
rect 263939 298392 263967 298420
rect 264001 298392 264029 298420
rect 264063 298392 264091 298420
rect 263877 290147 263905 290175
rect 263939 290147 263967 290175
rect 264001 290147 264029 290175
rect 264063 290147 264091 290175
rect 263877 290085 263905 290113
rect 263939 290085 263967 290113
rect 264001 290085 264029 290113
rect 264063 290085 264091 290113
rect 263877 290023 263905 290051
rect 263939 290023 263967 290051
rect 264001 290023 264029 290051
rect 264063 290023 264091 290051
rect 263877 289961 263905 289989
rect 263939 289961 263967 289989
rect 264001 289961 264029 289989
rect 264063 289961 264091 289989
rect 263877 281147 263905 281175
rect 263939 281147 263967 281175
rect 264001 281147 264029 281175
rect 264063 281147 264091 281175
rect 263877 281085 263905 281113
rect 263939 281085 263967 281113
rect 264001 281085 264029 281113
rect 264063 281085 264091 281113
rect 263877 281023 263905 281051
rect 263939 281023 263967 281051
rect 264001 281023 264029 281051
rect 264063 281023 264091 281051
rect 263877 280961 263905 280989
rect 263939 280961 263967 280989
rect 264001 280961 264029 280989
rect 264063 280961 264091 280989
rect 263877 272147 263905 272175
rect 263939 272147 263967 272175
rect 264001 272147 264029 272175
rect 264063 272147 264091 272175
rect 263877 272085 263905 272113
rect 263939 272085 263967 272113
rect 264001 272085 264029 272113
rect 264063 272085 264091 272113
rect 263877 272023 263905 272051
rect 263939 272023 263967 272051
rect 264001 272023 264029 272051
rect 264063 272023 264091 272051
rect 263877 271961 263905 271989
rect 263939 271961 263967 271989
rect 264001 271961 264029 271989
rect 264063 271961 264091 271989
rect 263877 263147 263905 263175
rect 263939 263147 263967 263175
rect 264001 263147 264029 263175
rect 264063 263147 264091 263175
rect 263877 263085 263905 263113
rect 263939 263085 263967 263113
rect 264001 263085 264029 263113
rect 264063 263085 264091 263113
rect 263877 263023 263905 263051
rect 263939 263023 263967 263051
rect 264001 263023 264029 263051
rect 264063 263023 264091 263051
rect 263877 262961 263905 262989
rect 263939 262961 263967 262989
rect 264001 262961 264029 262989
rect 264063 262961 264091 262989
rect 263877 254147 263905 254175
rect 263939 254147 263967 254175
rect 264001 254147 264029 254175
rect 264063 254147 264091 254175
rect 263877 254085 263905 254113
rect 263939 254085 263967 254113
rect 264001 254085 264029 254113
rect 264063 254085 264091 254113
rect 263877 254023 263905 254051
rect 263939 254023 263967 254051
rect 264001 254023 264029 254051
rect 264063 254023 264091 254051
rect 263877 253961 263905 253989
rect 263939 253961 263967 253989
rect 264001 253961 264029 253989
rect 264063 253961 264091 253989
rect 263877 245147 263905 245175
rect 263939 245147 263967 245175
rect 264001 245147 264029 245175
rect 264063 245147 264091 245175
rect 263877 245085 263905 245113
rect 263939 245085 263967 245113
rect 264001 245085 264029 245113
rect 264063 245085 264091 245113
rect 263877 245023 263905 245051
rect 263939 245023 263967 245051
rect 264001 245023 264029 245051
rect 264063 245023 264091 245051
rect 263877 244961 263905 244989
rect 263939 244961 263967 244989
rect 264001 244961 264029 244989
rect 264063 244961 264091 244989
rect 263877 236147 263905 236175
rect 263939 236147 263967 236175
rect 264001 236147 264029 236175
rect 264063 236147 264091 236175
rect 263877 236085 263905 236113
rect 263939 236085 263967 236113
rect 264001 236085 264029 236113
rect 264063 236085 264091 236113
rect 263877 236023 263905 236051
rect 263939 236023 263967 236051
rect 264001 236023 264029 236051
rect 264063 236023 264091 236051
rect 263877 235961 263905 235989
rect 263939 235961 263967 235989
rect 264001 235961 264029 235989
rect 264063 235961 264091 235989
rect 263877 227147 263905 227175
rect 263939 227147 263967 227175
rect 264001 227147 264029 227175
rect 264063 227147 264091 227175
rect 263877 227085 263905 227113
rect 263939 227085 263967 227113
rect 264001 227085 264029 227113
rect 264063 227085 264091 227113
rect 263877 227023 263905 227051
rect 263939 227023 263967 227051
rect 264001 227023 264029 227051
rect 264063 227023 264091 227051
rect 263877 226961 263905 226989
rect 263939 226961 263967 226989
rect 264001 226961 264029 226989
rect 264063 226961 264091 226989
rect 263877 218147 263905 218175
rect 263939 218147 263967 218175
rect 264001 218147 264029 218175
rect 264063 218147 264091 218175
rect 263877 218085 263905 218113
rect 263939 218085 263967 218113
rect 264001 218085 264029 218113
rect 264063 218085 264091 218113
rect 263877 218023 263905 218051
rect 263939 218023 263967 218051
rect 264001 218023 264029 218051
rect 264063 218023 264091 218051
rect 263877 217961 263905 217989
rect 263939 217961 263967 217989
rect 264001 217961 264029 217989
rect 264063 217961 264091 217989
rect 263877 209147 263905 209175
rect 263939 209147 263967 209175
rect 264001 209147 264029 209175
rect 264063 209147 264091 209175
rect 263877 209085 263905 209113
rect 263939 209085 263967 209113
rect 264001 209085 264029 209113
rect 264063 209085 264091 209113
rect 263877 209023 263905 209051
rect 263939 209023 263967 209051
rect 264001 209023 264029 209051
rect 264063 209023 264091 209051
rect 263877 208961 263905 208989
rect 263939 208961 263967 208989
rect 264001 208961 264029 208989
rect 264063 208961 264091 208989
rect 263877 200147 263905 200175
rect 263939 200147 263967 200175
rect 264001 200147 264029 200175
rect 264063 200147 264091 200175
rect 263877 200085 263905 200113
rect 263939 200085 263967 200113
rect 264001 200085 264029 200113
rect 264063 200085 264091 200113
rect 263877 200023 263905 200051
rect 263939 200023 263967 200051
rect 264001 200023 264029 200051
rect 264063 200023 264091 200051
rect 263877 199961 263905 199989
rect 263939 199961 263967 199989
rect 264001 199961 264029 199989
rect 264063 199961 264091 199989
rect 263877 191147 263905 191175
rect 263939 191147 263967 191175
rect 264001 191147 264029 191175
rect 264063 191147 264091 191175
rect 263877 191085 263905 191113
rect 263939 191085 263967 191113
rect 264001 191085 264029 191113
rect 264063 191085 264091 191113
rect 263877 191023 263905 191051
rect 263939 191023 263967 191051
rect 264001 191023 264029 191051
rect 264063 191023 264091 191051
rect 263877 190961 263905 190989
rect 263939 190961 263967 190989
rect 264001 190961 264029 190989
rect 264063 190961 264091 190989
rect 235017 185147 235045 185175
rect 235079 185147 235107 185175
rect 235141 185147 235169 185175
rect 235203 185147 235231 185175
rect 235017 185085 235045 185113
rect 235079 185085 235107 185113
rect 235141 185085 235169 185113
rect 235203 185085 235231 185113
rect 235017 185023 235045 185051
rect 235079 185023 235107 185051
rect 235141 185023 235169 185051
rect 235203 185023 235231 185051
rect 235017 184961 235045 184989
rect 235079 184961 235107 184989
rect 235141 184961 235169 184989
rect 235203 184961 235231 184989
rect 244939 185147 244967 185175
rect 245001 185147 245029 185175
rect 244939 185085 244967 185113
rect 245001 185085 245029 185113
rect 244939 185023 244967 185051
rect 245001 185023 245029 185051
rect 244939 184961 244967 184989
rect 245001 184961 245029 184989
rect 237259 182147 237287 182175
rect 237321 182147 237349 182175
rect 237259 182085 237287 182113
rect 237321 182085 237349 182113
rect 237259 182023 237287 182051
rect 237321 182023 237349 182051
rect 237259 181961 237287 181989
rect 237321 181961 237349 181989
rect 252619 182147 252647 182175
rect 252681 182147 252709 182175
rect 252619 182085 252647 182113
rect 252681 182085 252709 182113
rect 252619 182023 252647 182051
rect 252681 182023 252709 182051
rect 252619 181961 252647 181989
rect 252681 181961 252709 181989
rect 263877 182147 263905 182175
rect 263939 182147 263967 182175
rect 264001 182147 264029 182175
rect 264063 182147 264091 182175
rect 263877 182085 263905 182113
rect 263939 182085 263967 182113
rect 264001 182085 264029 182113
rect 264063 182085 264091 182113
rect 263877 182023 263905 182051
rect 263939 182023 263967 182051
rect 264001 182023 264029 182051
rect 264063 182023 264091 182051
rect 263877 181961 263905 181989
rect 263939 181961 263967 181989
rect 264001 181961 264029 181989
rect 264063 181961 264091 181989
rect 235017 176147 235045 176175
rect 235079 176147 235107 176175
rect 235141 176147 235169 176175
rect 235203 176147 235231 176175
rect 235017 176085 235045 176113
rect 235079 176085 235107 176113
rect 235141 176085 235169 176113
rect 235203 176085 235231 176113
rect 235017 176023 235045 176051
rect 235079 176023 235107 176051
rect 235141 176023 235169 176051
rect 235203 176023 235231 176051
rect 235017 175961 235045 175989
rect 235079 175961 235107 175989
rect 235141 175961 235169 175989
rect 235203 175961 235231 175989
rect 244939 176147 244967 176175
rect 245001 176147 245029 176175
rect 244939 176085 244967 176113
rect 245001 176085 245029 176113
rect 244939 176023 244967 176051
rect 245001 176023 245029 176051
rect 244939 175961 244967 175989
rect 245001 175961 245029 175989
rect 237259 173147 237287 173175
rect 237321 173147 237349 173175
rect 237259 173085 237287 173113
rect 237321 173085 237349 173113
rect 237259 173023 237287 173051
rect 237321 173023 237349 173051
rect 237259 172961 237287 172989
rect 237321 172961 237349 172989
rect 252619 173147 252647 173175
rect 252681 173147 252709 173175
rect 252619 173085 252647 173113
rect 252681 173085 252709 173113
rect 252619 173023 252647 173051
rect 252681 173023 252709 173051
rect 252619 172961 252647 172989
rect 252681 172961 252709 172989
rect 263877 173147 263905 173175
rect 263939 173147 263967 173175
rect 264001 173147 264029 173175
rect 264063 173147 264091 173175
rect 263877 173085 263905 173113
rect 263939 173085 263967 173113
rect 264001 173085 264029 173113
rect 264063 173085 264091 173113
rect 263877 173023 263905 173051
rect 263939 173023 263967 173051
rect 264001 173023 264029 173051
rect 264063 173023 264091 173051
rect 263877 172961 263905 172989
rect 263939 172961 263967 172989
rect 264001 172961 264029 172989
rect 264063 172961 264091 172989
rect 235017 167147 235045 167175
rect 235079 167147 235107 167175
rect 235141 167147 235169 167175
rect 235203 167147 235231 167175
rect 235017 167085 235045 167113
rect 235079 167085 235107 167113
rect 235141 167085 235169 167113
rect 235203 167085 235231 167113
rect 235017 167023 235045 167051
rect 235079 167023 235107 167051
rect 235141 167023 235169 167051
rect 235203 167023 235231 167051
rect 235017 166961 235045 166989
rect 235079 166961 235107 166989
rect 235141 166961 235169 166989
rect 235203 166961 235231 166989
rect 248517 164147 248545 164175
rect 248579 164147 248607 164175
rect 248641 164147 248669 164175
rect 248703 164147 248731 164175
rect 248517 164085 248545 164113
rect 248579 164085 248607 164113
rect 248641 164085 248669 164113
rect 248703 164085 248731 164113
rect 248517 164023 248545 164051
rect 248579 164023 248607 164051
rect 248641 164023 248669 164051
rect 248703 164023 248731 164051
rect 248517 163961 248545 163989
rect 248579 163961 248607 163989
rect 248641 163961 248669 163989
rect 248703 163961 248731 163989
rect 235017 158147 235045 158175
rect 235079 158147 235107 158175
rect 235141 158147 235169 158175
rect 235203 158147 235231 158175
rect 235017 158085 235045 158113
rect 235079 158085 235107 158113
rect 235141 158085 235169 158113
rect 235203 158085 235231 158113
rect 235017 158023 235045 158051
rect 235079 158023 235107 158051
rect 235141 158023 235169 158051
rect 235203 158023 235231 158051
rect 235017 157961 235045 157989
rect 235079 157961 235107 157989
rect 235141 157961 235169 157989
rect 235203 157961 235231 157989
rect 239619 158147 239647 158175
rect 239681 158147 239709 158175
rect 239619 158085 239647 158113
rect 239681 158085 239709 158113
rect 239619 158023 239647 158051
rect 239681 158023 239709 158051
rect 239619 157961 239647 157989
rect 239681 157961 239709 157989
rect 247299 155147 247327 155175
rect 247361 155147 247389 155175
rect 247299 155085 247327 155113
rect 247361 155085 247389 155113
rect 247299 155023 247327 155051
rect 247361 155023 247389 155051
rect 247299 154961 247327 154989
rect 247361 154961 247389 154989
rect 248517 155147 248545 155175
rect 248579 155147 248607 155175
rect 248641 155147 248669 155175
rect 248703 155147 248731 155175
rect 248517 155085 248545 155113
rect 248579 155085 248607 155113
rect 248641 155085 248669 155113
rect 248703 155085 248731 155113
rect 248517 155023 248545 155051
rect 248579 155023 248607 155051
rect 248641 155023 248669 155051
rect 248703 155023 248731 155051
rect 248517 154961 248545 154989
rect 248579 154961 248607 154989
rect 248641 154961 248669 154989
rect 248703 154961 248731 154989
rect 235017 149147 235045 149175
rect 235079 149147 235107 149175
rect 235141 149147 235169 149175
rect 235203 149147 235231 149175
rect 235017 149085 235045 149113
rect 235079 149085 235107 149113
rect 235141 149085 235169 149113
rect 235203 149085 235231 149113
rect 235017 149023 235045 149051
rect 235079 149023 235107 149051
rect 235141 149023 235169 149051
rect 235203 149023 235231 149051
rect 235017 148961 235045 148989
rect 235079 148961 235107 148989
rect 235141 148961 235169 148989
rect 235203 148961 235231 148989
rect 239619 149147 239647 149175
rect 239681 149147 239709 149175
rect 239619 149085 239647 149113
rect 239681 149085 239709 149113
rect 239619 149023 239647 149051
rect 239681 149023 239709 149051
rect 239619 148961 239647 148989
rect 239681 148961 239709 148989
rect 247299 146147 247327 146175
rect 247361 146147 247389 146175
rect 247299 146085 247327 146113
rect 247361 146085 247389 146113
rect 247299 146023 247327 146051
rect 247361 146023 247389 146051
rect 247299 145961 247327 145989
rect 247361 145961 247389 145989
rect 248517 146147 248545 146175
rect 248579 146147 248607 146175
rect 248641 146147 248669 146175
rect 248703 146147 248731 146175
rect 248517 146085 248545 146113
rect 248579 146085 248607 146113
rect 248641 146085 248669 146113
rect 248703 146085 248731 146113
rect 248517 146023 248545 146051
rect 248579 146023 248607 146051
rect 248641 146023 248669 146051
rect 248703 146023 248731 146051
rect 248517 145961 248545 145989
rect 248579 145961 248607 145989
rect 248641 145961 248669 145989
rect 248703 145961 248731 145989
rect 235017 140147 235045 140175
rect 235079 140147 235107 140175
rect 235141 140147 235169 140175
rect 235203 140147 235231 140175
rect 235017 140085 235045 140113
rect 235079 140085 235107 140113
rect 235141 140085 235169 140113
rect 235203 140085 235231 140113
rect 235017 140023 235045 140051
rect 235079 140023 235107 140051
rect 235141 140023 235169 140051
rect 235203 140023 235231 140051
rect 235017 139961 235045 139989
rect 235079 139961 235107 139989
rect 235141 139961 235169 139989
rect 235203 139961 235231 139989
rect 239619 140147 239647 140175
rect 239681 140147 239709 140175
rect 239619 140085 239647 140113
rect 239681 140085 239709 140113
rect 239619 140023 239647 140051
rect 239681 140023 239709 140051
rect 239619 139961 239647 139989
rect 239681 139961 239709 139989
rect 247299 137147 247327 137175
rect 247361 137147 247389 137175
rect 247299 137085 247327 137113
rect 247361 137085 247389 137113
rect 247299 137023 247327 137051
rect 247361 137023 247389 137051
rect 247299 136961 247327 136989
rect 247361 136961 247389 136989
rect 248517 137147 248545 137175
rect 248579 137147 248607 137175
rect 248641 137147 248669 137175
rect 248703 137147 248731 137175
rect 248517 137085 248545 137113
rect 248579 137085 248607 137113
rect 248641 137085 248669 137113
rect 248703 137085 248731 137113
rect 248517 137023 248545 137051
rect 248579 137023 248607 137051
rect 248641 137023 248669 137051
rect 248703 137023 248731 137051
rect 248517 136961 248545 136989
rect 248579 136961 248607 136989
rect 248641 136961 248669 136989
rect 248703 136961 248731 136989
rect 235017 131147 235045 131175
rect 235079 131147 235107 131175
rect 235141 131147 235169 131175
rect 235203 131147 235231 131175
rect 235017 131085 235045 131113
rect 235079 131085 235107 131113
rect 235141 131085 235169 131113
rect 235203 131085 235231 131113
rect 235017 131023 235045 131051
rect 235079 131023 235107 131051
rect 235141 131023 235169 131051
rect 235203 131023 235231 131051
rect 235017 130961 235045 130989
rect 235079 130961 235107 130989
rect 235141 130961 235169 130989
rect 235203 130961 235231 130989
rect 248517 128147 248545 128175
rect 248579 128147 248607 128175
rect 248641 128147 248669 128175
rect 248703 128147 248731 128175
rect 248517 128085 248545 128113
rect 248579 128085 248607 128113
rect 248641 128085 248669 128113
rect 248703 128085 248731 128113
rect 248517 128023 248545 128051
rect 248579 128023 248607 128051
rect 248641 128023 248669 128051
rect 248703 128023 248731 128051
rect 248517 127961 248545 127989
rect 248579 127961 248607 127989
rect 248641 127961 248669 127989
rect 248703 127961 248731 127989
rect 250377 167147 250405 167175
rect 250439 167147 250467 167175
rect 250501 167147 250529 167175
rect 250563 167147 250591 167175
rect 250377 167085 250405 167113
rect 250439 167085 250467 167113
rect 250501 167085 250529 167113
rect 250563 167085 250591 167113
rect 250377 167023 250405 167051
rect 250439 167023 250467 167051
rect 250501 167023 250529 167051
rect 250563 167023 250591 167051
rect 250377 166961 250405 166989
rect 250439 166961 250467 166989
rect 250501 166961 250529 166989
rect 250563 166961 250591 166989
rect 263877 164147 263905 164175
rect 263939 164147 263967 164175
rect 264001 164147 264029 164175
rect 264063 164147 264091 164175
rect 263877 164085 263905 164113
rect 263939 164085 263967 164113
rect 264001 164085 264029 164113
rect 264063 164085 264091 164113
rect 263877 164023 263905 164051
rect 263939 164023 263967 164051
rect 264001 164023 264029 164051
rect 264063 164023 264091 164051
rect 263877 163961 263905 163989
rect 263939 163961 263967 163989
rect 264001 163961 264029 163989
rect 264063 163961 264091 163989
rect 250377 158147 250405 158175
rect 250439 158147 250467 158175
rect 250501 158147 250529 158175
rect 250563 158147 250591 158175
rect 250377 158085 250405 158113
rect 250439 158085 250467 158113
rect 250501 158085 250529 158113
rect 250563 158085 250591 158113
rect 250377 158023 250405 158051
rect 250439 158023 250467 158051
rect 250501 158023 250529 158051
rect 250563 158023 250591 158051
rect 250377 157961 250405 157989
rect 250439 157961 250467 157989
rect 250501 157961 250529 157989
rect 250563 157961 250591 157989
rect 254979 158147 255007 158175
rect 255041 158147 255069 158175
rect 254979 158085 255007 158113
rect 255041 158085 255069 158113
rect 254979 158023 255007 158051
rect 255041 158023 255069 158051
rect 254979 157961 255007 157989
rect 255041 157961 255069 157989
rect 262659 155147 262687 155175
rect 262721 155147 262749 155175
rect 262659 155085 262687 155113
rect 262721 155085 262749 155113
rect 262659 155023 262687 155051
rect 262721 155023 262749 155051
rect 262659 154961 262687 154989
rect 262721 154961 262749 154989
rect 263877 155147 263905 155175
rect 263939 155147 263967 155175
rect 264001 155147 264029 155175
rect 264063 155147 264091 155175
rect 263877 155085 263905 155113
rect 263939 155085 263967 155113
rect 264001 155085 264029 155113
rect 264063 155085 264091 155113
rect 263877 155023 263905 155051
rect 263939 155023 263967 155051
rect 264001 155023 264029 155051
rect 264063 155023 264091 155051
rect 263877 154961 263905 154989
rect 263939 154961 263967 154989
rect 264001 154961 264029 154989
rect 264063 154961 264091 154989
rect 250377 149147 250405 149175
rect 250439 149147 250467 149175
rect 250501 149147 250529 149175
rect 250563 149147 250591 149175
rect 250377 149085 250405 149113
rect 250439 149085 250467 149113
rect 250501 149085 250529 149113
rect 250563 149085 250591 149113
rect 250377 149023 250405 149051
rect 250439 149023 250467 149051
rect 250501 149023 250529 149051
rect 250563 149023 250591 149051
rect 250377 148961 250405 148989
rect 250439 148961 250467 148989
rect 250501 148961 250529 148989
rect 250563 148961 250591 148989
rect 254979 149147 255007 149175
rect 255041 149147 255069 149175
rect 254979 149085 255007 149113
rect 255041 149085 255069 149113
rect 254979 149023 255007 149051
rect 255041 149023 255069 149051
rect 254979 148961 255007 148989
rect 255041 148961 255069 148989
rect 262659 146147 262687 146175
rect 262721 146147 262749 146175
rect 262659 146085 262687 146113
rect 262721 146085 262749 146113
rect 262659 146023 262687 146051
rect 262721 146023 262749 146051
rect 262659 145961 262687 145989
rect 262721 145961 262749 145989
rect 263877 146147 263905 146175
rect 263939 146147 263967 146175
rect 264001 146147 264029 146175
rect 264063 146147 264091 146175
rect 263877 146085 263905 146113
rect 263939 146085 263967 146113
rect 264001 146085 264029 146113
rect 264063 146085 264091 146113
rect 263877 146023 263905 146051
rect 263939 146023 263967 146051
rect 264001 146023 264029 146051
rect 264063 146023 264091 146051
rect 263877 145961 263905 145989
rect 263939 145961 263967 145989
rect 264001 145961 264029 145989
rect 264063 145961 264091 145989
rect 250377 140147 250405 140175
rect 250439 140147 250467 140175
rect 250501 140147 250529 140175
rect 250563 140147 250591 140175
rect 250377 140085 250405 140113
rect 250439 140085 250467 140113
rect 250501 140085 250529 140113
rect 250563 140085 250591 140113
rect 250377 140023 250405 140051
rect 250439 140023 250467 140051
rect 250501 140023 250529 140051
rect 250563 140023 250591 140051
rect 250377 139961 250405 139989
rect 250439 139961 250467 139989
rect 250501 139961 250529 139989
rect 250563 139961 250591 139989
rect 254979 140147 255007 140175
rect 255041 140147 255069 140175
rect 254979 140085 255007 140113
rect 255041 140085 255069 140113
rect 254979 140023 255007 140051
rect 255041 140023 255069 140051
rect 254979 139961 255007 139989
rect 255041 139961 255069 139989
rect 262659 137147 262687 137175
rect 262721 137147 262749 137175
rect 262659 137085 262687 137113
rect 262721 137085 262749 137113
rect 262659 137023 262687 137051
rect 262721 137023 262749 137051
rect 262659 136961 262687 136989
rect 262721 136961 262749 136989
rect 263877 137147 263905 137175
rect 263939 137147 263967 137175
rect 264001 137147 264029 137175
rect 264063 137147 264091 137175
rect 263877 137085 263905 137113
rect 263939 137085 263967 137113
rect 264001 137085 264029 137113
rect 264063 137085 264091 137113
rect 263877 137023 263905 137051
rect 263939 137023 263967 137051
rect 264001 137023 264029 137051
rect 264063 137023 264091 137051
rect 263877 136961 263905 136989
rect 263939 136961 263967 136989
rect 264001 136961 264029 136989
rect 264063 136961 264091 136989
rect 250377 131147 250405 131175
rect 250439 131147 250467 131175
rect 250501 131147 250529 131175
rect 250563 131147 250591 131175
rect 250377 131085 250405 131113
rect 250439 131085 250467 131113
rect 250501 131085 250529 131113
rect 250563 131085 250591 131113
rect 250377 131023 250405 131051
rect 250439 131023 250467 131051
rect 250501 131023 250529 131051
rect 250563 131023 250591 131051
rect 250377 130961 250405 130989
rect 250439 130961 250467 130989
rect 250501 130961 250529 130989
rect 250563 130961 250591 130989
rect 263877 128147 263905 128175
rect 263939 128147 263967 128175
rect 264001 128147 264029 128175
rect 264063 128147 264091 128175
rect 263877 128085 263905 128113
rect 263939 128085 263967 128113
rect 264001 128085 264029 128113
rect 264063 128085 264091 128113
rect 263877 128023 263905 128051
rect 263939 128023 263967 128051
rect 264001 128023 264029 128051
rect 264063 128023 264091 128051
rect 263877 127961 263905 127989
rect 263939 127961 263967 127989
rect 264001 127961 264029 127989
rect 264063 127961 264091 127989
rect 265737 299058 265765 299086
rect 265799 299058 265827 299086
rect 265861 299058 265889 299086
rect 265923 299058 265951 299086
rect 265737 298996 265765 299024
rect 265799 298996 265827 299024
rect 265861 298996 265889 299024
rect 265923 298996 265951 299024
rect 265737 298934 265765 298962
rect 265799 298934 265827 298962
rect 265861 298934 265889 298962
rect 265923 298934 265951 298962
rect 265737 298872 265765 298900
rect 265799 298872 265827 298900
rect 265861 298872 265889 298900
rect 265923 298872 265951 298900
rect 279237 298578 279265 298606
rect 279299 298578 279327 298606
rect 279361 298578 279389 298606
rect 279423 298578 279451 298606
rect 279237 298516 279265 298544
rect 279299 298516 279327 298544
rect 279361 298516 279389 298544
rect 279423 298516 279451 298544
rect 279237 298454 279265 298482
rect 279299 298454 279327 298482
rect 279361 298454 279389 298482
rect 279423 298454 279451 298482
rect 279237 298392 279265 298420
rect 279299 298392 279327 298420
rect 279361 298392 279389 298420
rect 279423 298392 279451 298420
rect 265737 293147 265765 293175
rect 265799 293147 265827 293175
rect 265861 293147 265889 293175
rect 265923 293147 265951 293175
rect 265737 293085 265765 293113
rect 265799 293085 265827 293113
rect 265861 293085 265889 293113
rect 265923 293085 265951 293113
rect 265737 293023 265765 293051
rect 265799 293023 265827 293051
rect 265861 293023 265889 293051
rect 265923 293023 265951 293051
rect 265737 292961 265765 292989
rect 265799 292961 265827 292989
rect 265861 292961 265889 292989
rect 265923 292961 265951 292989
rect 265737 284147 265765 284175
rect 265799 284147 265827 284175
rect 265861 284147 265889 284175
rect 265923 284147 265951 284175
rect 265737 284085 265765 284113
rect 265799 284085 265827 284113
rect 265861 284085 265889 284113
rect 265923 284085 265951 284113
rect 265737 284023 265765 284051
rect 265799 284023 265827 284051
rect 265861 284023 265889 284051
rect 265923 284023 265951 284051
rect 265737 283961 265765 283989
rect 265799 283961 265827 283989
rect 265861 283961 265889 283989
rect 265923 283961 265951 283989
rect 265737 275147 265765 275175
rect 265799 275147 265827 275175
rect 265861 275147 265889 275175
rect 265923 275147 265951 275175
rect 265737 275085 265765 275113
rect 265799 275085 265827 275113
rect 265861 275085 265889 275113
rect 265923 275085 265951 275113
rect 265737 275023 265765 275051
rect 265799 275023 265827 275051
rect 265861 275023 265889 275051
rect 265923 275023 265951 275051
rect 265737 274961 265765 274989
rect 265799 274961 265827 274989
rect 265861 274961 265889 274989
rect 265923 274961 265951 274989
rect 265737 266147 265765 266175
rect 265799 266147 265827 266175
rect 265861 266147 265889 266175
rect 265923 266147 265951 266175
rect 265737 266085 265765 266113
rect 265799 266085 265827 266113
rect 265861 266085 265889 266113
rect 265923 266085 265951 266113
rect 265737 266023 265765 266051
rect 265799 266023 265827 266051
rect 265861 266023 265889 266051
rect 265923 266023 265951 266051
rect 265737 265961 265765 265989
rect 265799 265961 265827 265989
rect 265861 265961 265889 265989
rect 265923 265961 265951 265989
rect 265737 257147 265765 257175
rect 265799 257147 265827 257175
rect 265861 257147 265889 257175
rect 265923 257147 265951 257175
rect 265737 257085 265765 257113
rect 265799 257085 265827 257113
rect 265861 257085 265889 257113
rect 265923 257085 265951 257113
rect 265737 257023 265765 257051
rect 265799 257023 265827 257051
rect 265861 257023 265889 257051
rect 265923 257023 265951 257051
rect 265737 256961 265765 256989
rect 265799 256961 265827 256989
rect 265861 256961 265889 256989
rect 265923 256961 265951 256989
rect 265737 248147 265765 248175
rect 265799 248147 265827 248175
rect 265861 248147 265889 248175
rect 265923 248147 265951 248175
rect 265737 248085 265765 248113
rect 265799 248085 265827 248113
rect 265861 248085 265889 248113
rect 265923 248085 265951 248113
rect 265737 248023 265765 248051
rect 265799 248023 265827 248051
rect 265861 248023 265889 248051
rect 265923 248023 265951 248051
rect 265737 247961 265765 247989
rect 265799 247961 265827 247989
rect 265861 247961 265889 247989
rect 265923 247961 265951 247989
rect 265737 239147 265765 239175
rect 265799 239147 265827 239175
rect 265861 239147 265889 239175
rect 265923 239147 265951 239175
rect 265737 239085 265765 239113
rect 265799 239085 265827 239113
rect 265861 239085 265889 239113
rect 265923 239085 265951 239113
rect 265737 239023 265765 239051
rect 265799 239023 265827 239051
rect 265861 239023 265889 239051
rect 265923 239023 265951 239051
rect 265737 238961 265765 238989
rect 265799 238961 265827 238989
rect 265861 238961 265889 238989
rect 265923 238961 265951 238989
rect 265737 230147 265765 230175
rect 265799 230147 265827 230175
rect 265861 230147 265889 230175
rect 265923 230147 265951 230175
rect 265737 230085 265765 230113
rect 265799 230085 265827 230113
rect 265861 230085 265889 230113
rect 265923 230085 265951 230113
rect 265737 230023 265765 230051
rect 265799 230023 265827 230051
rect 265861 230023 265889 230051
rect 265923 230023 265951 230051
rect 265737 229961 265765 229989
rect 265799 229961 265827 229989
rect 265861 229961 265889 229989
rect 265923 229961 265951 229989
rect 265737 221147 265765 221175
rect 265799 221147 265827 221175
rect 265861 221147 265889 221175
rect 265923 221147 265951 221175
rect 265737 221085 265765 221113
rect 265799 221085 265827 221113
rect 265861 221085 265889 221113
rect 265923 221085 265951 221113
rect 265737 221023 265765 221051
rect 265799 221023 265827 221051
rect 265861 221023 265889 221051
rect 265923 221023 265951 221051
rect 265737 220961 265765 220989
rect 265799 220961 265827 220989
rect 265861 220961 265889 220989
rect 265923 220961 265951 220989
rect 265737 212147 265765 212175
rect 265799 212147 265827 212175
rect 265861 212147 265889 212175
rect 265923 212147 265951 212175
rect 265737 212085 265765 212113
rect 265799 212085 265827 212113
rect 265861 212085 265889 212113
rect 265923 212085 265951 212113
rect 265737 212023 265765 212051
rect 265799 212023 265827 212051
rect 265861 212023 265889 212051
rect 265923 212023 265951 212051
rect 265737 211961 265765 211989
rect 265799 211961 265827 211989
rect 265861 211961 265889 211989
rect 265923 211961 265951 211989
rect 265737 203147 265765 203175
rect 265799 203147 265827 203175
rect 265861 203147 265889 203175
rect 265923 203147 265951 203175
rect 265737 203085 265765 203113
rect 265799 203085 265827 203113
rect 265861 203085 265889 203113
rect 265923 203085 265951 203113
rect 265737 203023 265765 203051
rect 265799 203023 265827 203051
rect 265861 203023 265889 203051
rect 265923 203023 265951 203051
rect 265737 202961 265765 202989
rect 265799 202961 265827 202989
rect 265861 202961 265889 202989
rect 265923 202961 265951 202989
rect 265737 194147 265765 194175
rect 265799 194147 265827 194175
rect 265861 194147 265889 194175
rect 265923 194147 265951 194175
rect 265737 194085 265765 194113
rect 265799 194085 265827 194113
rect 265861 194085 265889 194113
rect 265923 194085 265951 194113
rect 265737 194023 265765 194051
rect 265799 194023 265827 194051
rect 265861 194023 265889 194051
rect 265923 194023 265951 194051
rect 265737 193961 265765 193989
rect 265799 193961 265827 193989
rect 265861 193961 265889 193989
rect 265923 193961 265951 193989
rect 265737 185147 265765 185175
rect 265799 185147 265827 185175
rect 265861 185147 265889 185175
rect 265923 185147 265951 185175
rect 265737 185085 265765 185113
rect 265799 185085 265827 185113
rect 265861 185085 265889 185113
rect 265923 185085 265951 185113
rect 265737 185023 265765 185051
rect 265799 185023 265827 185051
rect 265861 185023 265889 185051
rect 265923 185023 265951 185051
rect 265737 184961 265765 184989
rect 265799 184961 265827 184989
rect 265861 184961 265889 184989
rect 265923 184961 265951 184989
rect 265737 176147 265765 176175
rect 265799 176147 265827 176175
rect 265861 176147 265889 176175
rect 265923 176147 265951 176175
rect 265737 176085 265765 176113
rect 265799 176085 265827 176113
rect 265861 176085 265889 176113
rect 265923 176085 265951 176113
rect 265737 176023 265765 176051
rect 265799 176023 265827 176051
rect 265861 176023 265889 176051
rect 265923 176023 265951 176051
rect 265737 175961 265765 175989
rect 265799 175961 265827 175989
rect 265861 175961 265889 175989
rect 265923 175961 265951 175989
rect 265737 167147 265765 167175
rect 265799 167147 265827 167175
rect 265861 167147 265889 167175
rect 265923 167147 265951 167175
rect 265737 167085 265765 167113
rect 265799 167085 265827 167113
rect 265861 167085 265889 167113
rect 265923 167085 265951 167113
rect 265737 167023 265765 167051
rect 265799 167023 265827 167051
rect 265861 167023 265889 167051
rect 265923 167023 265951 167051
rect 265737 166961 265765 166989
rect 265799 166961 265827 166989
rect 265861 166961 265889 166989
rect 265923 166961 265951 166989
rect 265737 158147 265765 158175
rect 265799 158147 265827 158175
rect 265861 158147 265889 158175
rect 265923 158147 265951 158175
rect 265737 158085 265765 158113
rect 265799 158085 265827 158113
rect 265861 158085 265889 158113
rect 265923 158085 265951 158113
rect 265737 158023 265765 158051
rect 265799 158023 265827 158051
rect 265861 158023 265889 158051
rect 265923 158023 265951 158051
rect 265737 157961 265765 157989
rect 265799 157961 265827 157989
rect 265861 157961 265889 157989
rect 265923 157961 265951 157989
rect 265737 149147 265765 149175
rect 265799 149147 265827 149175
rect 265861 149147 265889 149175
rect 265923 149147 265951 149175
rect 265737 149085 265765 149113
rect 265799 149085 265827 149113
rect 265861 149085 265889 149113
rect 265923 149085 265951 149113
rect 265737 149023 265765 149051
rect 265799 149023 265827 149051
rect 265861 149023 265889 149051
rect 265923 149023 265951 149051
rect 265737 148961 265765 148989
rect 265799 148961 265827 148989
rect 265861 148961 265889 148989
rect 265923 148961 265951 148989
rect 279237 290147 279265 290175
rect 279299 290147 279327 290175
rect 279361 290147 279389 290175
rect 279423 290147 279451 290175
rect 279237 290085 279265 290113
rect 279299 290085 279327 290113
rect 279361 290085 279389 290113
rect 279423 290085 279451 290113
rect 279237 290023 279265 290051
rect 279299 290023 279327 290051
rect 279361 290023 279389 290051
rect 279423 290023 279451 290051
rect 279237 289961 279265 289989
rect 279299 289961 279327 289989
rect 279361 289961 279389 289989
rect 279423 289961 279451 289989
rect 279237 281147 279265 281175
rect 279299 281147 279327 281175
rect 279361 281147 279389 281175
rect 279423 281147 279451 281175
rect 279237 281085 279265 281113
rect 279299 281085 279327 281113
rect 279361 281085 279389 281113
rect 279423 281085 279451 281113
rect 279237 281023 279265 281051
rect 279299 281023 279327 281051
rect 279361 281023 279389 281051
rect 279423 281023 279451 281051
rect 279237 280961 279265 280989
rect 279299 280961 279327 280989
rect 279361 280961 279389 280989
rect 279423 280961 279451 280989
rect 279237 272147 279265 272175
rect 279299 272147 279327 272175
rect 279361 272147 279389 272175
rect 279423 272147 279451 272175
rect 279237 272085 279265 272113
rect 279299 272085 279327 272113
rect 279361 272085 279389 272113
rect 279423 272085 279451 272113
rect 279237 272023 279265 272051
rect 279299 272023 279327 272051
rect 279361 272023 279389 272051
rect 279423 272023 279451 272051
rect 279237 271961 279265 271989
rect 279299 271961 279327 271989
rect 279361 271961 279389 271989
rect 279423 271961 279451 271989
rect 279237 263147 279265 263175
rect 279299 263147 279327 263175
rect 279361 263147 279389 263175
rect 279423 263147 279451 263175
rect 279237 263085 279265 263113
rect 279299 263085 279327 263113
rect 279361 263085 279389 263113
rect 279423 263085 279451 263113
rect 279237 263023 279265 263051
rect 279299 263023 279327 263051
rect 279361 263023 279389 263051
rect 279423 263023 279451 263051
rect 279237 262961 279265 262989
rect 279299 262961 279327 262989
rect 279361 262961 279389 262989
rect 279423 262961 279451 262989
rect 279237 254147 279265 254175
rect 279299 254147 279327 254175
rect 279361 254147 279389 254175
rect 279423 254147 279451 254175
rect 279237 254085 279265 254113
rect 279299 254085 279327 254113
rect 279361 254085 279389 254113
rect 279423 254085 279451 254113
rect 279237 254023 279265 254051
rect 279299 254023 279327 254051
rect 279361 254023 279389 254051
rect 279423 254023 279451 254051
rect 279237 253961 279265 253989
rect 279299 253961 279327 253989
rect 279361 253961 279389 253989
rect 279423 253961 279451 253989
rect 279237 245147 279265 245175
rect 279299 245147 279327 245175
rect 279361 245147 279389 245175
rect 279423 245147 279451 245175
rect 279237 245085 279265 245113
rect 279299 245085 279327 245113
rect 279361 245085 279389 245113
rect 279423 245085 279451 245113
rect 279237 245023 279265 245051
rect 279299 245023 279327 245051
rect 279361 245023 279389 245051
rect 279423 245023 279451 245051
rect 279237 244961 279265 244989
rect 279299 244961 279327 244989
rect 279361 244961 279389 244989
rect 279423 244961 279451 244989
rect 279237 236147 279265 236175
rect 279299 236147 279327 236175
rect 279361 236147 279389 236175
rect 279423 236147 279451 236175
rect 279237 236085 279265 236113
rect 279299 236085 279327 236113
rect 279361 236085 279389 236113
rect 279423 236085 279451 236113
rect 279237 236023 279265 236051
rect 279299 236023 279327 236051
rect 279361 236023 279389 236051
rect 279423 236023 279451 236051
rect 279237 235961 279265 235989
rect 279299 235961 279327 235989
rect 279361 235961 279389 235989
rect 279423 235961 279451 235989
rect 279237 227147 279265 227175
rect 279299 227147 279327 227175
rect 279361 227147 279389 227175
rect 279423 227147 279451 227175
rect 279237 227085 279265 227113
rect 279299 227085 279327 227113
rect 279361 227085 279389 227113
rect 279423 227085 279451 227113
rect 279237 227023 279265 227051
rect 279299 227023 279327 227051
rect 279361 227023 279389 227051
rect 279423 227023 279451 227051
rect 279237 226961 279265 226989
rect 279299 226961 279327 226989
rect 279361 226961 279389 226989
rect 279423 226961 279451 226989
rect 279237 218147 279265 218175
rect 279299 218147 279327 218175
rect 279361 218147 279389 218175
rect 279423 218147 279451 218175
rect 279237 218085 279265 218113
rect 279299 218085 279327 218113
rect 279361 218085 279389 218113
rect 279423 218085 279451 218113
rect 279237 218023 279265 218051
rect 279299 218023 279327 218051
rect 279361 218023 279389 218051
rect 279423 218023 279451 218051
rect 279237 217961 279265 217989
rect 279299 217961 279327 217989
rect 279361 217961 279389 217989
rect 279423 217961 279451 217989
rect 279237 209147 279265 209175
rect 279299 209147 279327 209175
rect 279361 209147 279389 209175
rect 279423 209147 279451 209175
rect 279237 209085 279265 209113
rect 279299 209085 279327 209113
rect 279361 209085 279389 209113
rect 279423 209085 279451 209113
rect 279237 209023 279265 209051
rect 279299 209023 279327 209051
rect 279361 209023 279389 209051
rect 279423 209023 279451 209051
rect 279237 208961 279265 208989
rect 279299 208961 279327 208989
rect 279361 208961 279389 208989
rect 279423 208961 279451 208989
rect 279237 200147 279265 200175
rect 279299 200147 279327 200175
rect 279361 200147 279389 200175
rect 279423 200147 279451 200175
rect 279237 200085 279265 200113
rect 279299 200085 279327 200113
rect 279361 200085 279389 200113
rect 279423 200085 279451 200113
rect 279237 200023 279265 200051
rect 279299 200023 279327 200051
rect 279361 200023 279389 200051
rect 279423 200023 279451 200051
rect 279237 199961 279265 199989
rect 279299 199961 279327 199989
rect 279361 199961 279389 199989
rect 279423 199961 279451 199989
rect 279237 191147 279265 191175
rect 279299 191147 279327 191175
rect 279361 191147 279389 191175
rect 279423 191147 279451 191175
rect 279237 191085 279265 191113
rect 279299 191085 279327 191113
rect 279361 191085 279389 191113
rect 279423 191085 279451 191113
rect 279237 191023 279265 191051
rect 279299 191023 279327 191051
rect 279361 191023 279389 191051
rect 279423 191023 279451 191051
rect 279237 190961 279265 190989
rect 279299 190961 279327 190989
rect 279361 190961 279389 190989
rect 279423 190961 279451 190989
rect 279237 182147 279265 182175
rect 279299 182147 279327 182175
rect 279361 182147 279389 182175
rect 279423 182147 279451 182175
rect 279237 182085 279265 182113
rect 279299 182085 279327 182113
rect 279361 182085 279389 182113
rect 279423 182085 279451 182113
rect 279237 182023 279265 182051
rect 279299 182023 279327 182051
rect 279361 182023 279389 182051
rect 279423 182023 279451 182051
rect 279237 181961 279265 181989
rect 279299 181961 279327 181989
rect 279361 181961 279389 181989
rect 279423 181961 279451 181989
rect 279237 173147 279265 173175
rect 279299 173147 279327 173175
rect 279361 173147 279389 173175
rect 279423 173147 279451 173175
rect 279237 173085 279265 173113
rect 279299 173085 279327 173113
rect 279361 173085 279389 173113
rect 279423 173085 279451 173113
rect 279237 173023 279265 173051
rect 279299 173023 279327 173051
rect 279361 173023 279389 173051
rect 279423 173023 279451 173051
rect 279237 172961 279265 172989
rect 279299 172961 279327 172989
rect 279361 172961 279389 172989
rect 279423 172961 279451 172989
rect 279237 164147 279265 164175
rect 279299 164147 279327 164175
rect 279361 164147 279389 164175
rect 279423 164147 279451 164175
rect 279237 164085 279265 164113
rect 279299 164085 279327 164113
rect 279361 164085 279389 164113
rect 279423 164085 279451 164113
rect 279237 164023 279265 164051
rect 279299 164023 279327 164051
rect 279361 164023 279389 164051
rect 279423 164023 279451 164051
rect 279237 163961 279265 163989
rect 279299 163961 279327 163989
rect 279361 163961 279389 163989
rect 279423 163961 279451 163989
rect 279237 155147 279265 155175
rect 279299 155147 279327 155175
rect 279361 155147 279389 155175
rect 279423 155147 279451 155175
rect 279237 155085 279265 155113
rect 279299 155085 279327 155113
rect 279361 155085 279389 155113
rect 279423 155085 279451 155113
rect 279237 155023 279265 155051
rect 279299 155023 279327 155051
rect 279361 155023 279389 155051
rect 279423 155023 279451 155051
rect 279237 154961 279265 154989
rect 279299 154961 279327 154989
rect 279361 154961 279389 154989
rect 279423 154961 279451 154989
rect 265737 140147 265765 140175
rect 265799 140147 265827 140175
rect 265861 140147 265889 140175
rect 265923 140147 265951 140175
rect 265737 140085 265765 140113
rect 265799 140085 265827 140113
rect 265861 140085 265889 140113
rect 265923 140085 265951 140113
rect 265737 140023 265765 140051
rect 265799 140023 265827 140051
rect 265861 140023 265889 140051
rect 265923 140023 265951 140051
rect 265737 139961 265765 139989
rect 265799 139961 265827 139989
rect 265861 139961 265889 139989
rect 265923 139961 265951 139989
rect 265737 131147 265765 131175
rect 265799 131147 265827 131175
rect 265861 131147 265889 131175
rect 265923 131147 265951 131175
rect 265737 131085 265765 131113
rect 265799 131085 265827 131113
rect 265861 131085 265889 131113
rect 265923 131085 265951 131113
rect 265737 131023 265765 131051
rect 265799 131023 265827 131051
rect 265861 131023 265889 131051
rect 265923 131023 265951 131051
rect 265737 130961 265765 130989
rect 265799 130961 265827 130989
rect 265861 130961 265889 130989
rect 265923 130961 265951 130989
rect 279237 146147 279265 146175
rect 279299 146147 279327 146175
rect 279361 146147 279389 146175
rect 279423 146147 279451 146175
rect 279237 146085 279265 146113
rect 279299 146085 279327 146113
rect 279361 146085 279389 146113
rect 279423 146085 279451 146113
rect 158217 122147 158245 122175
rect 158279 122147 158307 122175
rect 158341 122147 158369 122175
rect 158403 122147 158431 122175
rect 158217 122085 158245 122113
rect 158279 122085 158307 122113
rect 158341 122085 158369 122113
rect 158403 122085 158431 122113
rect 158217 122023 158245 122051
rect 158279 122023 158307 122051
rect 158341 122023 158369 122051
rect 158403 122023 158431 122051
rect 158217 121961 158245 121989
rect 158279 121961 158307 121989
rect 158341 121961 158369 121989
rect 158403 121961 158431 121989
rect 169939 122147 169967 122175
rect 170001 122147 170029 122175
rect 169939 122085 169967 122113
rect 170001 122085 170029 122113
rect 169939 122023 169967 122051
rect 170001 122023 170029 122051
rect 169939 121961 169967 121989
rect 170001 121961 170029 121989
rect 185299 122147 185327 122175
rect 185361 122147 185389 122175
rect 185299 122085 185327 122113
rect 185361 122085 185389 122113
rect 185299 122023 185327 122051
rect 185361 122023 185389 122051
rect 185299 121961 185327 121989
rect 185361 121961 185389 121989
rect 200659 122147 200687 122175
rect 200721 122147 200749 122175
rect 200659 122085 200687 122113
rect 200721 122085 200749 122113
rect 200659 122023 200687 122051
rect 200721 122023 200749 122051
rect 200659 121961 200687 121989
rect 200721 121961 200749 121989
rect 216019 122147 216047 122175
rect 216081 122147 216109 122175
rect 216019 122085 216047 122113
rect 216081 122085 216109 122113
rect 216019 122023 216047 122051
rect 216081 122023 216109 122051
rect 216019 121961 216047 121989
rect 216081 121961 216109 121989
rect 231379 122147 231407 122175
rect 231441 122147 231469 122175
rect 231379 122085 231407 122113
rect 231441 122085 231469 122113
rect 231379 122023 231407 122051
rect 231441 122023 231469 122051
rect 231379 121961 231407 121989
rect 231441 121961 231469 121989
rect 246739 122147 246767 122175
rect 246801 122147 246829 122175
rect 246739 122085 246767 122113
rect 246801 122085 246829 122113
rect 246739 122023 246767 122051
rect 246801 122023 246829 122051
rect 246739 121961 246767 121989
rect 246801 121961 246829 121989
rect 262099 122147 262127 122175
rect 262161 122147 262189 122175
rect 262099 122085 262127 122113
rect 262161 122085 262189 122113
rect 262099 122023 262127 122051
rect 262161 122023 262189 122051
rect 262099 121961 262127 121989
rect 262161 121961 262189 121989
rect 162259 119147 162287 119175
rect 162321 119147 162349 119175
rect 162259 119085 162287 119113
rect 162321 119085 162349 119113
rect 162259 119023 162287 119051
rect 162321 119023 162349 119051
rect 162259 118961 162287 118989
rect 162321 118961 162349 118989
rect 177619 119147 177647 119175
rect 177681 119147 177709 119175
rect 177619 119085 177647 119113
rect 177681 119085 177709 119113
rect 177619 119023 177647 119051
rect 177681 119023 177709 119051
rect 177619 118961 177647 118989
rect 177681 118961 177709 118989
rect 192979 119147 193007 119175
rect 193041 119147 193069 119175
rect 192979 119085 193007 119113
rect 193041 119085 193069 119113
rect 192979 119023 193007 119051
rect 193041 119023 193069 119051
rect 192979 118961 193007 118989
rect 193041 118961 193069 118989
rect 208339 119147 208367 119175
rect 208401 119147 208429 119175
rect 208339 119085 208367 119113
rect 208401 119085 208429 119113
rect 208339 119023 208367 119051
rect 208401 119023 208429 119051
rect 208339 118961 208367 118989
rect 208401 118961 208429 118989
rect 223699 119147 223727 119175
rect 223761 119147 223789 119175
rect 223699 119085 223727 119113
rect 223761 119085 223789 119113
rect 223699 119023 223727 119051
rect 223761 119023 223789 119051
rect 223699 118961 223727 118989
rect 223761 118961 223789 118989
rect 239059 119147 239087 119175
rect 239121 119147 239149 119175
rect 239059 119085 239087 119113
rect 239121 119085 239149 119113
rect 239059 119023 239087 119051
rect 239121 119023 239149 119051
rect 239059 118961 239087 118989
rect 239121 118961 239149 118989
rect 254419 119147 254447 119175
rect 254481 119147 254509 119175
rect 254419 119085 254447 119113
rect 254481 119085 254509 119113
rect 254419 119023 254447 119051
rect 254481 119023 254509 119051
rect 254419 118961 254447 118989
rect 254481 118961 254509 118989
rect 269779 119147 269807 119175
rect 269841 119147 269869 119175
rect 269779 119085 269807 119113
rect 269841 119085 269869 119113
rect 269779 119023 269807 119051
rect 269841 119023 269869 119051
rect 269779 118961 269807 118989
rect 269841 118961 269869 118989
rect 158217 113147 158245 113175
rect 158279 113147 158307 113175
rect 158341 113147 158369 113175
rect 158403 113147 158431 113175
rect 158217 113085 158245 113113
rect 158279 113085 158307 113113
rect 158341 113085 158369 113113
rect 158403 113085 158431 113113
rect 158217 113023 158245 113051
rect 158279 113023 158307 113051
rect 158341 113023 158369 113051
rect 158403 113023 158431 113051
rect 158217 112961 158245 112989
rect 158279 112961 158307 112989
rect 158341 112961 158369 112989
rect 158403 112961 158431 112989
rect 169939 113147 169967 113175
rect 170001 113147 170029 113175
rect 169939 113085 169967 113113
rect 170001 113085 170029 113113
rect 169939 113023 169967 113051
rect 170001 113023 170029 113051
rect 169939 112961 169967 112989
rect 170001 112961 170029 112989
rect 185299 113147 185327 113175
rect 185361 113147 185389 113175
rect 185299 113085 185327 113113
rect 185361 113085 185389 113113
rect 185299 113023 185327 113051
rect 185361 113023 185389 113051
rect 185299 112961 185327 112989
rect 185361 112961 185389 112989
rect 200659 113147 200687 113175
rect 200721 113147 200749 113175
rect 200659 113085 200687 113113
rect 200721 113085 200749 113113
rect 200659 113023 200687 113051
rect 200721 113023 200749 113051
rect 200659 112961 200687 112989
rect 200721 112961 200749 112989
rect 216019 113147 216047 113175
rect 216081 113147 216109 113175
rect 216019 113085 216047 113113
rect 216081 113085 216109 113113
rect 216019 113023 216047 113051
rect 216081 113023 216109 113051
rect 216019 112961 216047 112989
rect 216081 112961 216109 112989
rect 231379 113147 231407 113175
rect 231441 113147 231469 113175
rect 231379 113085 231407 113113
rect 231441 113085 231469 113113
rect 231379 113023 231407 113051
rect 231441 113023 231469 113051
rect 231379 112961 231407 112989
rect 231441 112961 231469 112989
rect 246739 113147 246767 113175
rect 246801 113147 246829 113175
rect 246739 113085 246767 113113
rect 246801 113085 246829 113113
rect 246739 113023 246767 113051
rect 246801 113023 246829 113051
rect 246739 112961 246767 112989
rect 246801 112961 246829 112989
rect 262099 113147 262127 113175
rect 262161 113147 262189 113175
rect 262099 113085 262127 113113
rect 262161 113085 262189 113113
rect 262099 113023 262127 113051
rect 262161 113023 262189 113051
rect 262099 112961 262127 112989
rect 262161 112961 262189 112989
rect 162259 110147 162287 110175
rect 162321 110147 162349 110175
rect 162259 110085 162287 110113
rect 162321 110085 162349 110113
rect 162259 110023 162287 110051
rect 162321 110023 162349 110051
rect 162259 109961 162287 109989
rect 162321 109961 162349 109989
rect 177619 110147 177647 110175
rect 177681 110147 177709 110175
rect 177619 110085 177647 110113
rect 177681 110085 177709 110113
rect 177619 110023 177647 110051
rect 177681 110023 177709 110051
rect 177619 109961 177647 109989
rect 177681 109961 177709 109989
rect 192979 110147 193007 110175
rect 193041 110147 193069 110175
rect 192979 110085 193007 110113
rect 193041 110085 193069 110113
rect 192979 110023 193007 110051
rect 193041 110023 193069 110051
rect 192979 109961 193007 109989
rect 193041 109961 193069 109989
rect 208339 110147 208367 110175
rect 208401 110147 208429 110175
rect 208339 110085 208367 110113
rect 208401 110085 208429 110113
rect 208339 110023 208367 110051
rect 208401 110023 208429 110051
rect 208339 109961 208367 109989
rect 208401 109961 208429 109989
rect 223699 110147 223727 110175
rect 223761 110147 223789 110175
rect 223699 110085 223727 110113
rect 223761 110085 223789 110113
rect 223699 110023 223727 110051
rect 223761 110023 223789 110051
rect 223699 109961 223727 109989
rect 223761 109961 223789 109989
rect 239059 110147 239087 110175
rect 239121 110147 239149 110175
rect 239059 110085 239087 110113
rect 239121 110085 239149 110113
rect 239059 110023 239087 110051
rect 239121 110023 239149 110051
rect 239059 109961 239087 109989
rect 239121 109961 239149 109989
rect 254419 110147 254447 110175
rect 254481 110147 254509 110175
rect 254419 110085 254447 110113
rect 254481 110085 254509 110113
rect 254419 110023 254447 110051
rect 254481 110023 254509 110051
rect 254419 109961 254447 109989
rect 254481 109961 254509 109989
rect 269779 110147 269807 110175
rect 269841 110147 269869 110175
rect 269779 110085 269807 110113
rect 269841 110085 269869 110113
rect 269779 110023 269807 110051
rect 269841 110023 269869 110051
rect 269779 109961 269807 109989
rect 269841 109961 269869 109989
rect 158217 104147 158245 104175
rect 158279 104147 158307 104175
rect 158341 104147 158369 104175
rect 158403 104147 158431 104175
rect 158217 104085 158245 104113
rect 158279 104085 158307 104113
rect 158341 104085 158369 104113
rect 158403 104085 158431 104113
rect 158217 104023 158245 104051
rect 158279 104023 158307 104051
rect 158341 104023 158369 104051
rect 158403 104023 158431 104051
rect 158217 103961 158245 103989
rect 158279 103961 158307 103989
rect 158341 103961 158369 103989
rect 158403 103961 158431 103989
rect 169939 104147 169967 104175
rect 170001 104147 170029 104175
rect 169939 104085 169967 104113
rect 170001 104085 170029 104113
rect 169939 104023 169967 104051
rect 170001 104023 170029 104051
rect 169939 103961 169967 103989
rect 170001 103961 170029 103989
rect 185299 104147 185327 104175
rect 185361 104147 185389 104175
rect 185299 104085 185327 104113
rect 185361 104085 185389 104113
rect 185299 104023 185327 104051
rect 185361 104023 185389 104051
rect 185299 103961 185327 103989
rect 185361 103961 185389 103989
rect 200659 104147 200687 104175
rect 200721 104147 200749 104175
rect 200659 104085 200687 104113
rect 200721 104085 200749 104113
rect 200659 104023 200687 104051
rect 200721 104023 200749 104051
rect 200659 103961 200687 103989
rect 200721 103961 200749 103989
rect 216019 104147 216047 104175
rect 216081 104147 216109 104175
rect 216019 104085 216047 104113
rect 216081 104085 216109 104113
rect 216019 104023 216047 104051
rect 216081 104023 216109 104051
rect 216019 103961 216047 103989
rect 216081 103961 216109 103989
rect 231379 104147 231407 104175
rect 231441 104147 231469 104175
rect 231379 104085 231407 104113
rect 231441 104085 231469 104113
rect 231379 104023 231407 104051
rect 231441 104023 231469 104051
rect 231379 103961 231407 103989
rect 231441 103961 231469 103989
rect 246739 104147 246767 104175
rect 246801 104147 246829 104175
rect 246739 104085 246767 104113
rect 246801 104085 246829 104113
rect 246739 104023 246767 104051
rect 246801 104023 246829 104051
rect 246739 103961 246767 103989
rect 246801 103961 246829 103989
rect 262099 104147 262127 104175
rect 262161 104147 262189 104175
rect 262099 104085 262127 104113
rect 262161 104085 262189 104113
rect 262099 104023 262127 104051
rect 262161 104023 262189 104051
rect 262099 103961 262127 103989
rect 262161 103961 262189 103989
rect 162259 101147 162287 101175
rect 162321 101147 162349 101175
rect 162259 101085 162287 101113
rect 162321 101085 162349 101113
rect 162259 101023 162287 101051
rect 162321 101023 162349 101051
rect 162259 100961 162287 100989
rect 162321 100961 162349 100989
rect 177619 101147 177647 101175
rect 177681 101147 177709 101175
rect 177619 101085 177647 101113
rect 177681 101085 177709 101113
rect 177619 101023 177647 101051
rect 177681 101023 177709 101051
rect 177619 100961 177647 100989
rect 177681 100961 177709 100989
rect 192979 101147 193007 101175
rect 193041 101147 193069 101175
rect 192979 101085 193007 101113
rect 193041 101085 193069 101113
rect 192979 101023 193007 101051
rect 193041 101023 193069 101051
rect 192979 100961 193007 100989
rect 193041 100961 193069 100989
rect 208339 101147 208367 101175
rect 208401 101147 208429 101175
rect 208339 101085 208367 101113
rect 208401 101085 208429 101113
rect 208339 101023 208367 101051
rect 208401 101023 208429 101051
rect 208339 100961 208367 100989
rect 208401 100961 208429 100989
rect 223699 101147 223727 101175
rect 223761 101147 223789 101175
rect 223699 101085 223727 101113
rect 223761 101085 223789 101113
rect 223699 101023 223727 101051
rect 223761 101023 223789 101051
rect 223699 100961 223727 100989
rect 223761 100961 223789 100989
rect 239059 101147 239087 101175
rect 239121 101147 239149 101175
rect 239059 101085 239087 101113
rect 239121 101085 239149 101113
rect 239059 101023 239087 101051
rect 239121 101023 239149 101051
rect 239059 100961 239087 100989
rect 239121 100961 239149 100989
rect 254419 101147 254447 101175
rect 254481 101147 254509 101175
rect 254419 101085 254447 101113
rect 254481 101085 254509 101113
rect 254419 101023 254447 101051
rect 254481 101023 254509 101051
rect 254419 100961 254447 100989
rect 254481 100961 254509 100989
rect 269779 101147 269807 101175
rect 269841 101147 269869 101175
rect 269779 101085 269807 101113
rect 269841 101085 269869 101113
rect 269779 101023 269807 101051
rect 269841 101023 269869 101051
rect 269779 100961 269807 100989
rect 269841 100961 269869 100989
rect 158217 95147 158245 95175
rect 158279 95147 158307 95175
rect 158341 95147 158369 95175
rect 158403 95147 158431 95175
rect 158217 95085 158245 95113
rect 158279 95085 158307 95113
rect 158341 95085 158369 95113
rect 158403 95085 158431 95113
rect 158217 95023 158245 95051
rect 158279 95023 158307 95051
rect 158341 95023 158369 95051
rect 158403 95023 158431 95051
rect 158217 94961 158245 94989
rect 158279 94961 158307 94989
rect 158341 94961 158369 94989
rect 158403 94961 158431 94989
rect 169939 95147 169967 95175
rect 170001 95147 170029 95175
rect 169939 95085 169967 95113
rect 170001 95085 170029 95113
rect 169939 95023 169967 95051
rect 170001 95023 170029 95051
rect 169939 94961 169967 94989
rect 170001 94961 170029 94989
rect 185299 95147 185327 95175
rect 185361 95147 185389 95175
rect 185299 95085 185327 95113
rect 185361 95085 185389 95113
rect 185299 95023 185327 95051
rect 185361 95023 185389 95051
rect 185299 94961 185327 94989
rect 185361 94961 185389 94989
rect 200659 95147 200687 95175
rect 200721 95147 200749 95175
rect 200659 95085 200687 95113
rect 200721 95085 200749 95113
rect 200659 95023 200687 95051
rect 200721 95023 200749 95051
rect 200659 94961 200687 94989
rect 200721 94961 200749 94989
rect 216019 95147 216047 95175
rect 216081 95147 216109 95175
rect 216019 95085 216047 95113
rect 216081 95085 216109 95113
rect 216019 95023 216047 95051
rect 216081 95023 216109 95051
rect 216019 94961 216047 94989
rect 216081 94961 216109 94989
rect 231379 95147 231407 95175
rect 231441 95147 231469 95175
rect 231379 95085 231407 95113
rect 231441 95085 231469 95113
rect 231379 95023 231407 95051
rect 231441 95023 231469 95051
rect 231379 94961 231407 94989
rect 231441 94961 231469 94989
rect 246739 95147 246767 95175
rect 246801 95147 246829 95175
rect 246739 95085 246767 95113
rect 246801 95085 246829 95113
rect 246739 95023 246767 95051
rect 246801 95023 246829 95051
rect 246739 94961 246767 94989
rect 246801 94961 246829 94989
rect 262099 95147 262127 95175
rect 262161 95147 262189 95175
rect 262099 95085 262127 95113
rect 262161 95085 262189 95113
rect 262099 95023 262127 95051
rect 262161 95023 262189 95051
rect 262099 94961 262127 94989
rect 262161 94961 262189 94989
rect 162259 92147 162287 92175
rect 162321 92147 162349 92175
rect 162259 92085 162287 92113
rect 162321 92085 162349 92113
rect 162259 92023 162287 92051
rect 162321 92023 162349 92051
rect 162259 91961 162287 91989
rect 162321 91961 162349 91989
rect 177619 92147 177647 92175
rect 177681 92147 177709 92175
rect 177619 92085 177647 92113
rect 177681 92085 177709 92113
rect 177619 92023 177647 92051
rect 177681 92023 177709 92051
rect 177619 91961 177647 91989
rect 177681 91961 177709 91989
rect 192979 92147 193007 92175
rect 193041 92147 193069 92175
rect 192979 92085 193007 92113
rect 193041 92085 193069 92113
rect 192979 92023 193007 92051
rect 193041 92023 193069 92051
rect 192979 91961 193007 91989
rect 193041 91961 193069 91989
rect 208339 92147 208367 92175
rect 208401 92147 208429 92175
rect 208339 92085 208367 92113
rect 208401 92085 208429 92113
rect 208339 92023 208367 92051
rect 208401 92023 208429 92051
rect 208339 91961 208367 91989
rect 208401 91961 208429 91989
rect 223699 92147 223727 92175
rect 223761 92147 223789 92175
rect 223699 92085 223727 92113
rect 223761 92085 223789 92113
rect 223699 92023 223727 92051
rect 223761 92023 223789 92051
rect 223699 91961 223727 91989
rect 223761 91961 223789 91989
rect 239059 92147 239087 92175
rect 239121 92147 239149 92175
rect 239059 92085 239087 92113
rect 239121 92085 239149 92113
rect 239059 92023 239087 92051
rect 239121 92023 239149 92051
rect 239059 91961 239087 91989
rect 239121 91961 239149 91989
rect 254419 92147 254447 92175
rect 254481 92147 254509 92175
rect 254419 92085 254447 92113
rect 254481 92085 254509 92113
rect 254419 92023 254447 92051
rect 254481 92023 254509 92051
rect 254419 91961 254447 91989
rect 254481 91961 254509 91989
rect 269779 92147 269807 92175
rect 269841 92147 269869 92175
rect 269779 92085 269807 92113
rect 269841 92085 269869 92113
rect 269779 92023 269807 92051
rect 269841 92023 269869 92051
rect 269779 91961 269807 91989
rect 269841 91961 269869 91989
rect 158217 86147 158245 86175
rect 158279 86147 158307 86175
rect 158341 86147 158369 86175
rect 158403 86147 158431 86175
rect 158217 86085 158245 86113
rect 158279 86085 158307 86113
rect 158341 86085 158369 86113
rect 158403 86085 158431 86113
rect 158217 86023 158245 86051
rect 158279 86023 158307 86051
rect 158341 86023 158369 86051
rect 158403 86023 158431 86051
rect 158217 85961 158245 85989
rect 158279 85961 158307 85989
rect 158341 85961 158369 85989
rect 158403 85961 158431 85989
rect 169939 86147 169967 86175
rect 170001 86147 170029 86175
rect 169939 86085 169967 86113
rect 170001 86085 170029 86113
rect 169939 86023 169967 86051
rect 170001 86023 170029 86051
rect 169939 85961 169967 85989
rect 170001 85961 170029 85989
rect 185299 86147 185327 86175
rect 185361 86147 185389 86175
rect 185299 86085 185327 86113
rect 185361 86085 185389 86113
rect 185299 86023 185327 86051
rect 185361 86023 185389 86051
rect 185299 85961 185327 85989
rect 185361 85961 185389 85989
rect 200659 86147 200687 86175
rect 200721 86147 200749 86175
rect 200659 86085 200687 86113
rect 200721 86085 200749 86113
rect 200659 86023 200687 86051
rect 200721 86023 200749 86051
rect 200659 85961 200687 85989
rect 200721 85961 200749 85989
rect 216019 86147 216047 86175
rect 216081 86147 216109 86175
rect 216019 86085 216047 86113
rect 216081 86085 216109 86113
rect 216019 86023 216047 86051
rect 216081 86023 216109 86051
rect 216019 85961 216047 85989
rect 216081 85961 216109 85989
rect 231379 86147 231407 86175
rect 231441 86147 231469 86175
rect 231379 86085 231407 86113
rect 231441 86085 231469 86113
rect 231379 86023 231407 86051
rect 231441 86023 231469 86051
rect 231379 85961 231407 85989
rect 231441 85961 231469 85989
rect 246739 86147 246767 86175
rect 246801 86147 246829 86175
rect 246739 86085 246767 86113
rect 246801 86085 246829 86113
rect 246739 86023 246767 86051
rect 246801 86023 246829 86051
rect 246739 85961 246767 85989
rect 246801 85961 246829 85989
rect 262099 86147 262127 86175
rect 262161 86147 262189 86175
rect 262099 86085 262127 86113
rect 262161 86085 262189 86113
rect 262099 86023 262127 86051
rect 262161 86023 262189 86051
rect 262099 85961 262127 85989
rect 262161 85961 262189 85989
rect 162259 83147 162287 83175
rect 162321 83147 162349 83175
rect 162259 83085 162287 83113
rect 162321 83085 162349 83113
rect 162259 83023 162287 83051
rect 162321 83023 162349 83051
rect 162259 82961 162287 82989
rect 162321 82961 162349 82989
rect 177619 83147 177647 83175
rect 177681 83147 177709 83175
rect 177619 83085 177647 83113
rect 177681 83085 177709 83113
rect 177619 83023 177647 83051
rect 177681 83023 177709 83051
rect 177619 82961 177647 82989
rect 177681 82961 177709 82989
rect 192979 83147 193007 83175
rect 193041 83147 193069 83175
rect 192979 83085 193007 83113
rect 193041 83085 193069 83113
rect 192979 83023 193007 83051
rect 193041 83023 193069 83051
rect 192979 82961 193007 82989
rect 193041 82961 193069 82989
rect 208339 83147 208367 83175
rect 208401 83147 208429 83175
rect 208339 83085 208367 83113
rect 208401 83085 208429 83113
rect 208339 83023 208367 83051
rect 208401 83023 208429 83051
rect 208339 82961 208367 82989
rect 208401 82961 208429 82989
rect 223699 83147 223727 83175
rect 223761 83147 223789 83175
rect 223699 83085 223727 83113
rect 223761 83085 223789 83113
rect 223699 83023 223727 83051
rect 223761 83023 223789 83051
rect 223699 82961 223727 82989
rect 223761 82961 223789 82989
rect 239059 83147 239087 83175
rect 239121 83147 239149 83175
rect 239059 83085 239087 83113
rect 239121 83085 239149 83113
rect 239059 83023 239087 83051
rect 239121 83023 239149 83051
rect 239059 82961 239087 82989
rect 239121 82961 239149 82989
rect 254419 83147 254447 83175
rect 254481 83147 254509 83175
rect 254419 83085 254447 83113
rect 254481 83085 254509 83113
rect 254419 83023 254447 83051
rect 254481 83023 254509 83051
rect 254419 82961 254447 82989
rect 254481 82961 254509 82989
rect 269779 83147 269807 83175
rect 269841 83147 269869 83175
rect 269779 83085 269807 83113
rect 269841 83085 269869 83113
rect 269779 83023 269807 83051
rect 269841 83023 269869 83051
rect 269779 82961 269807 82989
rect 269841 82961 269869 82989
rect 158217 77147 158245 77175
rect 158279 77147 158307 77175
rect 158341 77147 158369 77175
rect 158403 77147 158431 77175
rect 158217 77085 158245 77113
rect 158279 77085 158307 77113
rect 158341 77085 158369 77113
rect 158403 77085 158431 77113
rect 158217 77023 158245 77051
rect 158279 77023 158307 77051
rect 158341 77023 158369 77051
rect 158403 77023 158431 77051
rect 158217 76961 158245 76989
rect 158279 76961 158307 76989
rect 158341 76961 158369 76989
rect 158403 76961 158431 76989
rect 169939 77147 169967 77175
rect 170001 77147 170029 77175
rect 169939 77085 169967 77113
rect 170001 77085 170029 77113
rect 169939 77023 169967 77051
rect 170001 77023 170029 77051
rect 169939 76961 169967 76989
rect 170001 76961 170029 76989
rect 185299 77147 185327 77175
rect 185361 77147 185389 77175
rect 185299 77085 185327 77113
rect 185361 77085 185389 77113
rect 185299 77023 185327 77051
rect 185361 77023 185389 77051
rect 185299 76961 185327 76989
rect 185361 76961 185389 76989
rect 200659 77147 200687 77175
rect 200721 77147 200749 77175
rect 200659 77085 200687 77113
rect 200721 77085 200749 77113
rect 200659 77023 200687 77051
rect 200721 77023 200749 77051
rect 200659 76961 200687 76989
rect 200721 76961 200749 76989
rect 216019 77147 216047 77175
rect 216081 77147 216109 77175
rect 216019 77085 216047 77113
rect 216081 77085 216109 77113
rect 216019 77023 216047 77051
rect 216081 77023 216109 77051
rect 216019 76961 216047 76989
rect 216081 76961 216109 76989
rect 231379 77147 231407 77175
rect 231441 77147 231469 77175
rect 231379 77085 231407 77113
rect 231441 77085 231469 77113
rect 231379 77023 231407 77051
rect 231441 77023 231469 77051
rect 231379 76961 231407 76989
rect 231441 76961 231469 76989
rect 246739 77147 246767 77175
rect 246801 77147 246829 77175
rect 246739 77085 246767 77113
rect 246801 77085 246829 77113
rect 246739 77023 246767 77051
rect 246801 77023 246829 77051
rect 246739 76961 246767 76989
rect 246801 76961 246829 76989
rect 262099 77147 262127 77175
rect 262161 77147 262189 77175
rect 262099 77085 262127 77113
rect 262161 77085 262189 77113
rect 262099 77023 262127 77051
rect 262161 77023 262189 77051
rect 262099 76961 262127 76989
rect 262161 76961 262189 76989
rect 162259 74147 162287 74175
rect 162321 74147 162349 74175
rect 162259 74085 162287 74113
rect 162321 74085 162349 74113
rect 162259 74023 162287 74051
rect 162321 74023 162349 74051
rect 162259 73961 162287 73989
rect 162321 73961 162349 73989
rect 177619 74147 177647 74175
rect 177681 74147 177709 74175
rect 177619 74085 177647 74113
rect 177681 74085 177709 74113
rect 177619 74023 177647 74051
rect 177681 74023 177709 74051
rect 177619 73961 177647 73989
rect 177681 73961 177709 73989
rect 192979 74147 193007 74175
rect 193041 74147 193069 74175
rect 192979 74085 193007 74113
rect 193041 74085 193069 74113
rect 192979 74023 193007 74051
rect 193041 74023 193069 74051
rect 192979 73961 193007 73989
rect 193041 73961 193069 73989
rect 208339 74147 208367 74175
rect 208401 74147 208429 74175
rect 208339 74085 208367 74113
rect 208401 74085 208429 74113
rect 208339 74023 208367 74051
rect 208401 74023 208429 74051
rect 208339 73961 208367 73989
rect 208401 73961 208429 73989
rect 223699 74147 223727 74175
rect 223761 74147 223789 74175
rect 223699 74085 223727 74113
rect 223761 74085 223789 74113
rect 223699 74023 223727 74051
rect 223761 74023 223789 74051
rect 223699 73961 223727 73989
rect 223761 73961 223789 73989
rect 239059 74147 239087 74175
rect 239121 74147 239149 74175
rect 239059 74085 239087 74113
rect 239121 74085 239149 74113
rect 239059 74023 239087 74051
rect 239121 74023 239149 74051
rect 239059 73961 239087 73989
rect 239121 73961 239149 73989
rect 254419 74147 254447 74175
rect 254481 74147 254509 74175
rect 254419 74085 254447 74113
rect 254481 74085 254509 74113
rect 254419 74023 254447 74051
rect 254481 74023 254509 74051
rect 254419 73961 254447 73989
rect 254481 73961 254509 73989
rect 269779 74147 269807 74175
rect 269841 74147 269869 74175
rect 269779 74085 269807 74113
rect 269841 74085 269869 74113
rect 269779 74023 269807 74051
rect 269841 74023 269869 74051
rect 269779 73961 269807 73989
rect 269841 73961 269869 73989
rect 158217 68147 158245 68175
rect 158279 68147 158307 68175
rect 158341 68147 158369 68175
rect 158403 68147 158431 68175
rect 158217 68085 158245 68113
rect 158279 68085 158307 68113
rect 158341 68085 158369 68113
rect 158403 68085 158431 68113
rect 158217 68023 158245 68051
rect 158279 68023 158307 68051
rect 158341 68023 158369 68051
rect 158403 68023 158431 68051
rect 158217 67961 158245 67989
rect 158279 67961 158307 67989
rect 158341 67961 158369 67989
rect 158403 67961 158431 67989
rect 169939 68147 169967 68175
rect 170001 68147 170029 68175
rect 169939 68085 169967 68113
rect 170001 68085 170029 68113
rect 169939 68023 169967 68051
rect 170001 68023 170029 68051
rect 169939 67961 169967 67989
rect 170001 67961 170029 67989
rect 185299 68147 185327 68175
rect 185361 68147 185389 68175
rect 185299 68085 185327 68113
rect 185361 68085 185389 68113
rect 185299 68023 185327 68051
rect 185361 68023 185389 68051
rect 185299 67961 185327 67989
rect 185361 67961 185389 67989
rect 200659 68147 200687 68175
rect 200721 68147 200749 68175
rect 200659 68085 200687 68113
rect 200721 68085 200749 68113
rect 200659 68023 200687 68051
rect 200721 68023 200749 68051
rect 200659 67961 200687 67989
rect 200721 67961 200749 67989
rect 216019 68147 216047 68175
rect 216081 68147 216109 68175
rect 216019 68085 216047 68113
rect 216081 68085 216109 68113
rect 216019 68023 216047 68051
rect 216081 68023 216109 68051
rect 216019 67961 216047 67989
rect 216081 67961 216109 67989
rect 231379 68147 231407 68175
rect 231441 68147 231469 68175
rect 231379 68085 231407 68113
rect 231441 68085 231469 68113
rect 231379 68023 231407 68051
rect 231441 68023 231469 68051
rect 231379 67961 231407 67989
rect 231441 67961 231469 67989
rect 246739 68147 246767 68175
rect 246801 68147 246829 68175
rect 246739 68085 246767 68113
rect 246801 68085 246829 68113
rect 246739 68023 246767 68051
rect 246801 68023 246829 68051
rect 246739 67961 246767 67989
rect 246801 67961 246829 67989
rect 262099 68147 262127 68175
rect 262161 68147 262189 68175
rect 262099 68085 262127 68113
rect 262161 68085 262189 68113
rect 262099 68023 262127 68051
rect 262161 68023 262189 68051
rect 262099 67961 262127 67989
rect 262161 67961 262189 67989
rect 162259 65147 162287 65175
rect 162321 65147 162349 65175
rect 162259 65085 162287 65113
rect 162321 65085 162349 65113
rect 162259 65023 162287 65051
rect 162321 65023 162349 65051
rect 162259 64961 162287 64989
rect 162321 64961 162349 64989
rect 177619 65147 177647 65175
rect 177681 65147 177709 65175
rect 177619 65085 177647 65113
rect 177681 65085 177709 65113
rect 177619 65023 177647 65051
rect 177681 65023 177709 65051
rect 177619 64961 177647 64989
rect 177681 64961 177709 64989
rect 192979 65147 193007 65175
rect 193041 65147 193069 65175
rect 192979 65085 193007 65113
rect 193041 65085 193069 65113
rect 192979 65023 193007 65051
rect 193041 65023 193069 65051
rect 192979 64961 193007 64989
rect 193041 64961 193069 64989
rect 208339 65147 208367 65175
rect 208401 65147 208429 65175
rect 208339 65085 208367 65113
rect 208401 65085 208429 65113
rect 208339 65023 208367 65051
rect 208401 65023 208429 65051
rect 208339 64961 208367 64989
rect 208401 64961 208429 64989
rect 223699 65147 223727 65175
rect 223761 65147 223789 65175
rect 223699 65085 223727 65113
rect 223761 65085 223789 65113
rect 223699 65023 223727 65051
rect 223761 65023 223789 65051
rect 223699 64961 223727 64989
rect 223761 64961 223789 64989
rect 239059 65147 239087 65175
rect 239121 65147 239149 65175
rect 239059 65085 239087 65113
rect 239121 65085 239149 65113
rect 239059 65023 239087 65051
rect 239121 65023 239149 65051
rect 239059 64961 239087 64989
rect 239121 64961 239149 64989
rect 254419 65147 254447 65175
rect 254481 65147 254509 65175
rect 254419 65085 254447 65113
rect 254481 65085 254509 65113
rect 254419 65023 254447 65051
rect 254481 65023 254509 65051
rect 254419 64961 254447 64989
rect 254481 64961 254509 64989
rect 269779 65147 269807 65175
rect 269841 65147 269869 65175
rect 269779 65085 269807 65113
rect 269841 65085 269869 65113
rect 269779 65023 269807 65051
rect 269841 65023 269869 65051
rect 269779 64961 269807 64989
rect 269841 64961 269869 64989
rect 158217 59147 158245 59175
rect 158279 59147 158307 59175
rect 158341 59147 158369 59175
rect 158403 59147 158431 59175
rect 158217 59085 158245 59113
rect 158279 59085 158307 59113
rect 158341 59085 158369 59113
rect 158403 59085 158431 59113
rect 158217 59023 158245 59051
rect 158279 59023 158307 59051
rect 158341 59023 158369 59051
rect 158403 59023 158431 59051
rect 158217 58961 158245 58989
rect 158279 58961 158307 58989
rect 158341 58961 158369 58989
rect 158403 58961 158431 58989
rect 169939 59147 169967 59175
rect 170001 59147 170029 59175
rect 169939 59085 169967 59113
rect 170001 59085 170029 59113
rect 169939 59023 169967 59051
rect 170001 59023 170029 59051
rect 169939 58961 169967 58989
rect 170001 58961 170029 58989
rect 185299 59147 185327 59175
rect 185361 59147 185389 59175
rect 185299 59085 185327 59113
rect 185361 59085 185389 59113
rect 185299 59023 185327 59051
rect 185361 59023 185389 59051
rect 185299 58961 185327 58989
rect 185361 58961 185389 58989
rect 200659 59147 200687 59175
rect 200721 59147 200749 59175
rect 200659 59085 200687 59113
rect 200721 59085 200749 59113
rect 200659 59023 200687 59051
rect 200721 59023 200749 59051
rect 200659 58961 200687 58989
rect 200721 58961 200749 58989
rect 216019 59147 216047 59175
rect 216081 59147 216109 59175
rect 216019 59085 216047 59113
rect 216081 59085 216109 59113
rect 216019 59023 216047 59051
rect 216081 59023 216109 59051
rect 216019 58961 216047 58989
rect 216081 58961 216109 58989
rect 231379 59147 231407 59175
rect 231441 59147 231469 59175
rect 231379 59085 231407 59113
rect 231441 59085 231469 59113
rect 231379 59023 231407 59051
rect 231441 59023 231469 59051
rect 231379 58961 231407 58989
rect 231441 58961 231469 58989
rect 246739 59147 246767 59175
rect 246801 59147 246829 59175
rect 246739 59085 246767 59113
rect 246801 59085 246829 59113
rect 246739 59023 246767 59051
rect 246801 59023 246829 59051
rect 246739 58961 246767 58989
rect 246801 58961 246829 58989
rect 262099 59147 262127 59175
rect 262161 59147 262189 59175
rect 262099 59085 262127 59113
rect 262161 59085 262189 59113
rect 262099 59023 262127 59051
rect 262161 59023 262189 59051
rect 262099 58961 262127 58989
rect 262161 58961 262189 58989
rect 162259 56147 162287 56175
rect 162321 56147 162349 56175
rect 162259 56085 162287 56113
rect 162321 56085 162349 56113
rect 162259 56023 162287 56051
rect 162321 56023 162349 56051
rect 162259 55961 162287 55989
rect 162321 55961 162349 55989
rect 177619 56147 177647 56175
rect 177681 56147 177709 56175
rect 177619 56085 177647 56113
rect 177681 56085 177709 56113
rect 177619 56023 177647 56051
rect 177681 56023 177709 56051
rect 177619 55961 177647 55989
rect 177681 55961 177709 55989
rect 192979 56147 193007 56175
rect 193041 56147 193069 56175
rect 192979 56085 193007 56113
rect 193041 56085 193069 56113
rect 192979 56023 193007 56051
rect 193041 56023 193069 56051
rect 192979 55961 193007 55989
rect 193041 55961 193069 55989
rect 208339 56147 208367 56175
rect 208401 56147 208429 56175
rect 208339 56085 208367 56113
rect 208401 56085 208429 56113
rect 208339 56023 208367 56051
rect 208401 56023 208429 56051
rect 208339 55961 208367 55989
rect 208401 55961 208429 55989
rect 223699 56147 223727 56175
rect 223761 56147 223789 56175
rect 223699 56085 223727 56113
rect 223761 56085 223789 56113
rect 223699 56023 223727 56051
rect 223761 56023 223789 56051
rect 223699 55961 223727 55989
rect 223761 55961 223789 55989
rect 239059 56147 239087 56175
rect 239121 56147 239149 56175
rect 239059 56085 239087 56113
rect 239121 56085 239149 56113
rect 239059 56023 239087 56051
rect 239121 56023 239149 56051
rect 239059 55961 239087 55989
rect 239121 55961 239149 55989
rect 254419 56147 254447 56175
rect 254481 56147 254509 56175
rect 254419 56085 254447 56113
rect 254481 56085 254509 56113
rect 254419 56023 254447 56051
rect 254481 56023 254509 56051
rect 254419 55961 254447 55989
rect 254481 55961 254509 55989
rect 269779 56147 269807 56175
rect 269841 56147 269869 56175
rect 269779 56085 269807 56113
rect 269841 56085 269869 56113
rect 269779 56023 269807 56051
rect 269841 56023 269869 56051
rect 269779 55961 269807 55989
rect 269841 55961 269869 55989
rect 158217 50147 158245 50175
rect 158279 50147 158307 50175
rect 158341 50147 158369 50175
rect 158403 50147 158431 50175
rect 158217 50085 158245 50113
rect 158279 50085 158307 50113
rect 158341 50085 158369 50113
rect 158403 50085 158431 50113
rect 158217 50023 158245 50051
rect 158279 50023 158307 50051
rect 158341 50023 158369 50051
rect 158403 50023 158431 50051
rect 158217 49961 158245 49989
rect 158279 49961 158307 49989
rect 158341 49961 158369 49989
rect 158403 49961 158431 49989
rect 169939 50147 169967 50175
rect 170001 50147 170029 50175
rect 169939 50085 169967 50113
rect 170001 50085 170029 50113
rect 169939 50023 169967 50051
rect 170001 50023 170029 50051
rect 169939 49961 169967 49989
rect 170001 49961 170029 49989
rect 185299 50147 185327 50175
rect 185361 50147 185389 50175
rect 185299 50085 185327 50113
rect 185361 50085 185389 50113
rect 185299 50023 185327 50051
rect 185361 50023 185389 50051
rect 185299 49961 185327 49989
rect 185361 49961 185389 49989
rect 200659 50147 200687 50175
rect 200721 50147 200749 50175
rect 200659 50085 200687 50113
rect 200721 50085 200749 50113
rect 200659 50023 200687 50051
rect 200721 50023 200749 50051
rect 200659 49961 200687 49989
rect 200721 49961 200749 49989
rect 216019 50147 216047 50175
rect 216081 50147 216109 50175
rect 216019 50085 216047 50113
rect 216081 50085 216109 50113
rect 216019 50023 216047 50051
rect 216081 50023 216109 50051
rect 216019 49961 216047 49989
rect 216081 49961 216109 49989
rect 231379 50147 231407 50175
rect 231441 50147 231469 50175
rect 231379 50085 231407 50113
rect 231441 50085 231469 50113
rect 231379 50023 231407 50051
rect 231441 50023 231469 50051
rect 231379 49961 231407 49989
rect 231441 49961 231469 49989
rect 246739 50147 246767 50175
rect 246801 50147 246829 50175
rect 246739 50085 246767 50113
rect 246801 50085 246829 50113
rect 246739 50023 246767 50051
rect 246801 50023 246829 50051
rect 246739 49961 246767 49989
rect 246801 49961 246829 49989
rect 262099 50147 262127 50175
rect 262161 50147 262189 50175
rect 262099 50085 262127 50113
rect 262161 50085 262189 50113
rect 262099 50023 262127 50051
rect 262161 50023 262189 50051
rect 262099 49961 262127 49989
rect 262161 49961 262189 49989
rect 162259 47147 162287 47175
rect 162321 47147 162349 47175
rect 162259 47085 162287 47113
rect 162321 47085 162349 47113
rect 162259 47023 162287 47051
rect 162321 47023 162349 47051
rect 162259 46961 162287 46989
rect 162321 46961 162349 46989
rect 177619 47147 177647 47175
rect 177681 47147 177709 47175
rect 177619 47085 177647 47113
rect 177681 47085 177709 47113
rect 177619 47023 177647 47051
rect 177681 47023 177709 47051
rect 177619 46961 177647 46989
rect 177681 46961 177709 46989
rect 192979 47147 193007 47175
rect 193041 47147 193069 47175
rect 192979 47085 193007 47113
rect 193041 47085 193069 47113
rect 192979 47023 193007 47051
rect 193041 47023 193069 47051
rect 192979 46961 193007 46989
rect 193041 46961 193069 46989
rect 208339 47147 208367 47175
rect 208401 47147 208429 47175
rect 208339 47085 208367 47113
rect 208401 47085 208429 47113
rect 208339 47023 208367 47051
rect 208401 47023 208429 47051
rect 208339 46961 208367 46989
rect 208401 46961 208429 46989
rect 223699 47147 223727 47175
rect 223761 47147 223789 47175
rect 223699 47085 223727 47113
rect 223761 47085 223789 47113
rect 223699 47023 223727 47051
rect 223761 47023 223789 47051
rect 223699 46961 223727 46989
rect 223761 46961 223789 46989
rect 239059 47147 239087 47175
rect 239121 47147 239149 47175
rect 239059 47085 239087 47113
rect 239121 47085 239149 47113
rect 239059 47023 239087 47051
rect 239121 47023 239149 47051
rect 239059 46961 239087 46989
rect 239121 46961 239149 46989
rect 254419 47147 254447 47175
rect 254481 47147 254509 47175
rect 254419 47085 254447 47113
rect 254481 47085 254509 47113
rect 254419 47023 254447 47051
rect 254481 47023 254509 47051
rect 254419 46961 254447 46989
rect 254481 46961 254509 46989
rect 269779 47147 269807 47175
rect 269841 47147 269869 47175
rect 269779 47085 269807 47113
rect 269841 47085 269869 47113
rect 269779 47023 269807 47051
rect 269841 47023 269869 47051
rect 269779 46961 269807 46989
rect 269841 46961 269869 46989
rect 158217 41147 158245 41175
rect 158279 41147 158307 41175
rect 158341 41147 158369 41175
rect 158403 41147 158431 41175
rect 158217 41085 158245 41113
rect 158279 41085 158307 41113
rect 158341 41085 158369 41113
rect 158403 41085 158431 41113
rect 158217 41023 158245 41051
rect 158279 41023 158307 41051
rect 158341 41023 158369 41051
rect 158403 41023 158431 41051
rect 158217 40961 158245 40989
rect 158279 40961 158307 40989
rect 158341 40961 158369 40989
rect 158403 40961 158431 40989
rect 169939 41147 169967 41175
rect 170001 41147 170029 41175
rect 169939 41085 169967 41113
rect 170001 41085 170029 41113
rect 169939 41023 169967 41051
rect 170001 41023 170029 41051
rect 169939 40961 169967 40989
rect 170001 40961 170029 40989
rect 185299 41147 185327 41175
rect 185361 41147 185389 41175
rect 185299 41085 185327 41113
rect 185361 41085 185389 41113
rect 185299 41023 185327 41051
rect 185361 41023 185389 41051
rect 185299 40961 185327 40989
rect 185361 40961 185389 40989
rect 200659 41147 200687 41175
rect 200721 41147 200749 41175
rect 200659 41085 200687 41113
rect 200721 41085 200749 41113
rect 200659 41023 200687 41051
rect 200721 41023 200749 41051
rect 200659 40961 200687 40989
rect 200721 40961 200749 40989
rect 216019 41147 216047 41175
rect 216081 41147 216109 41175
rect 216019 41085 216047 41113
rect 216081 41085 216109 41113
rect 216019 41023 216047 41051
rect 216081 41023 216109 41051
rect 216019 40961 216047 40989
rect 216081 40961 216109 40989
rect 231379 41147 231407 41175
rect 231441 41147 231469 41175
rect 231379 41085 231407 41113
rect 231441 41085 231469 41113
rect 231379 41023 231407 41051
rect 231441 41023 231469 41051
rect 231379 40961 231407 40989
rect 231441 40961 231469 40989
rect 246739 41147 246767 41175
rect 246801 41147 246829 41175
rect 246739 41085 246767 41113
rect 246801 41085 246829 41113
rect 246739 41023 246767 41051
rect 246801 41023 246829 41051
rect 246739 40961 246767 40989
rect 246801 40961 246829 40989
rect 262099 41147 262127 41175
rect 262161 41147 262189 41175
rect 262099 41085 262127 41113
rect 262161 41085 262189 41113
rect 262099 41023 262127 41051
rect 262161 41023 262189 41051
rect 262099 40961 262127 40989
rect 262161 40961 262189 40989
rect 162259 38147 162287 38175
rect 162321 38147 162349 38175
rect 162259 38085 162287 38113
rect 162321 38085 162349 38113
rect 162259 38023 162287 38051
rect 162321 38023 162349 38051
rect 162259 37961 162287 37989
rect 162321 37961 162349 37989
rect 177619 38147 177647 38175
rect 177681 38147 177709 38175
rect 177619 38085 177647 38113
rect 177681 38085 177709 38113
rect 177619 38023 177647 38051
rect 177681 38023 177709 38051
rect 177619 37961 177647 37989
rect 177681 37961 177709 37989
rect 192979 38147 193007 38175
rect 193041 38147 193069 38175
rect 192979 38085 193007 38113
rect 193041 38085 193069 38113
rect 192979 38023 193007 38051
rect 193041 38023 193069 38051
rect 192979 37961 193007 37989
rect 193041 37961 193069 37989
rect 208339 38147 208367 38175
rect 208401 38147 208429 38175
rect 208339 38085 208367 38113
rect 208401 38085 208429 38113
rect 208339 38023 208367 38051
rect 208401 38023 208429 38051
rect 208339 37961 208367 37989
rect 208401 37961 208429 37989
rect 223699 38147 223727 38175
rect 223761 38147 223789 38175
rect 223699 38085 223727 38113
rect 223761 38085 223789 38113
rect 223699 38023 223727 38051
rect 223761 38023 223789 38051
rect 223699 37961 223727 37989
rect 223761 37961 223789 37989
rect 239059 38147 239087 38175
rect 239121 38147 239149 38175
rect 239059 38085 239087 38113
rect 239121 38085 239149 38113
rect 239059 38023 239087 38051
rect 239121 38023 239149 38051
rect 239059 37961 239087 37989
rect 239121 37961 239149 37989
rect 254419 38147 254447 38175
rect 254481 38147 254509 38175
rect 254419 38085 254447 38113
rect 254481 38085 254509 38113
rect 254419 38023 254447 38051
rect 254481 38023 254509 38051
rect 254419 37961 254447 37989
rect 254481 37961 254509 37989
rect 269779 38147 269807 38175
rect 269841 38147 269869 38175
rect 269779 38085 269807 38113
rect 269841 38085 269869 38113
rect 269779 38023 269807 38051
rect 269841 38023 269869 38051
rect 269779 37961 269807 37989
rect 269841 37961 269869 37989
rect 158217 32147 158245 32175
rect 158279 32147 158307 32175
rect 158341 32147 158369 32175
rect 158403 32147 158431 32175
rect 158217 32085 158245 32113
rect 158279 32085 158307 32113
rect 158341 32085 158369 32113
rect 158403 32085 158431 32113
rect 158217 32023 158245 32051
rect 158279 32023 158307 32051
rect 158341 32023 158369 32051
rect 158403 32023 158431 32051
rect 158217 31961 158245 31989
rect 158279 31961 158307 31989
rect 158341 31961 158369 31989
rect 158403 31961 158431 31989
rect 169939 32147 169967 32175
rect 170001 32147 170029 32175
rect 169939 32085 169967 32113
rect 170001 32085 170029 32113
rect 169939 32023 169967 32051
rect 170001 32023 170029 32051
rect 169939 31961 169967 31989
rect 170001 31961 170029 31989
rect 185299 32147 185327 32175
rect 185361 32147 185389 32175
rect 185299 32085 185327 32113
rect 185361 32085 185389 32113
rect 185299 32023 185327 32051
rect 185361 32023 185389 32051
rect 185299 31961 185327 31989
rect 185361 31961 185389 31989
rect 200659 32147 200687 32175
rect 200721 32147 200749 32175
rect 200659 32085 200687 32113
rect 200721 32085 200749 32113
rect 200659 32023 200687 32051
rect 200721 32023 200749 32051
rect 200659 31961 200687 31989
rect 200721 31961 200749 31989
rect 216019 32147 216047 32175
rect 216081 32147 216109 32175
rect 216019 32085 216047 32113
rect 216081 32085 216109 32113
rect 216019 32023 216047 32051
rect 216081 32023 216109 32051
rect 216019 31961 216047 31989
rect 216081 31961 216109 31989
rect 231379 32147 231407 32175
rect 231441 32147 231469 32175
rect 231379 32085 231407 32113
rect 231441 32085 231469 32113
rect 231379 32023 231407 32051
rect 231441 32023 231469 32051
rect 231379 31961 231407 31989
rect 231441 31961 231469 31989
rect 246739 32147 246767 32175
rect 246801 32147 246829 32175
rect 246739 32085 246767 32113
rect 246801 32085 246829 32113
rect 246739 32023 246767 32051
rect 246801 32023 246829 32051
rect 246739 31961 246767 31989
rect 246801 31961 246829 31989
rect 262099 32147 262127 32175
rect 262161 32147 262189 32175
rect 262099 32085 262127 32113
rect 262161 32085 262189 32113
rect 262099 32023 262127 32051
rect 262161 32023 262189 32051
rect 262099 31961 262127 31989
rect 262161 31961 262189 31989
rect 162259 29147 162287 29175
rect 162321 29147 162349 29175
rect 162259 29085 162287 29113
rect 162321 29085 162349 29113
rect 162259 29023 162287 29051
rect 162321 29023 162349 29051
rect 162259 28961 162287 28989
rect 162321 28961 162349 28989
rect 177619 29147 177647 29175
rect 177681 29147 177709 29175
rect 177619 29085 177647 29113
rect 177681 29085 177709 29113
rect 177619 29023 177647 29051
rect 177681 29023 177709 29051
rect 177619 28961 177647 28989
rect 177681 28961 177709 28989
rect 192979 29147 193007 29175
rect 193041 29147 193069 29175
rect 192979 29085 193007 29113
rect 193041 29085 193069 29113
rect 192979 29023 193007 29051
rect 193041 29023 193069 29051
rect 192979 28961 193007 28989
rect 193041 28961 193069 28989
rect 208339 29147 208367 29175
rect 208401 29147 208429 29175
rect 208339 29085 208367 29113
rect 208401 29085 208429 29113
rect 208339 29023 208367 29051
rect 208401 29023 208429 29051
rect 208339 28961 208367 28989
rect 208401 28961 208429 28989
rect 223699 29147 223727 29175
rect 223761 29147 223789 29175
rect 223699 29085 223727 29113
rect 223761 29085 223789 29113
rect 223699 29023 223727 29051
rect 223761 29023 223789 29051
rect 223699 28961 223727 28989
rect 223761 28961 223789 28989
rect 239059 29147 239087 29175
rect 239121 29147 239149 29175
rect 239059 29085 239087 29113
rect 239121 29085 239149 29113
rect 239059 29023 239087 29051
rect 239121 29023 239149 29051
rect 239059 28961 239087 28989
rect 239121 28961 239149 28989
rect 254419 29147 254447 29175
rect 254481 29147 254509 29175
rect 254419 29085 254447 29113
rect 254481 29085 254509 29113
rect 254419 29023 254447 29051
rect 254481 29023 254509 29051
rect 254419 28961 254447 28989
rect 254481 28961 254509 28989
rect 269779 29147 269807 29175
rect 269841 29147 269869 29175
rect 269779 29085 269807 29113
rect 269841 29085 269869 29113
rect 269779 29023 269807 29051
rect 269841 29023 269869 29051
rect 269779 28961 269807 28989
rect 269841 28961 269869 28989
rect 158217 23147 158245 23175
rect 158279 23147 158307 23175
rect 158341 23147 158369 23175
rect 158403 23147 158431 23175
rect 158217 23085 158245 23113
rect 158279 23085 158307 23113
rect 158341 23085 158369 23113
rect 158403 23085 158431 23113
rect 158217 23023 158245 23051
rect 158279 23023 158307 23051
rect 158341 23023 158369 23051
rect 158403 23023 158431 23051
rect 158217 22961 158245 22989
rect 158279 22961 158307 22989
rect 158341 22961 158369 22989
rect 158403 22961 158431 22989
rect 169939 23147 169967 23175
rect 170001 23147 170029 23175
rect 169939 23085 169967 23113
rect 170001 23085 170029 23113
rect 169939 23023 169967 23051
rect 170001 23023 170029 23051
rect 169939 22961 169967 22989
rect 170001 22961 170029 22989
rect 185299 23147 185327 23175
rect 185361 23147 185389 23175
rect 185299 23085 185327 23113
rect 185361 23085 185389 23113
rect 185299 23023 185327 23051
rect 185361 23023 185389 23051
rect 185299 22961 185327 22989
rect 185361 22961 185389 22989
rect 200659 23147 200687 23175
rect 200721 23147 200749 23175
rect 200659 23085 200687 23113
rect 200721 23085 200749 23113
rect 200659 23023 200687 23051
rect 200721 23023 200749 23051
rect 200659 22961 200687 22989
rect 200721 22961 200749 22989
rect 216019 23147 216047 23175
rect 216081 23147 216109 23175
rect 216019 23085 216047 23113
rect 216081 23085 216109 23113
rect 216019 23023 216047 23051
rect 216081 23023 216109 23051
rect 216019 22961 216047 22989
rect 216081 22961 216109 22989
rect 231379 23147 231407 23175
rect 231441 23147 231469 23175
rect 231379 23085 231407 23113
rect 231441 23085 231469 23113
rect 231379 23023 231407 23051
rect 231441 23023 231469 23051
rect 231379 22961 231407 22989
rect 231441 22961 231469 22989
rect 246739 23147 246767 23175
rect 246801 23147 246829 23175
rect 246739 23085 246767 23113
rect 246801 23085 246829 23113
rect 246739 23023 246767 23051
rect 246801 23023 246829 23051
rect 246739 22961 246767 22989
rect 246801 22961 246829 22989
rect 262099 23147 262127 23175
rect 262161 23147 262189 23175
rect 262099 23085 262127 23113
rect 262161 23085 262189 23113
rect 262099 23023 262127 23051
rect 262161 23023 262189 23051
rect 262099 22961 262127 22989
rect 262161 22961 262189 22989
rect 162259 20147 162287 20175
rect 162321 20147 162349 20175
rect 162259 20085 162287 20113
rect 162321 20085 162349 20113
rect 162259 20023 162287 20051
rect 162321 20023 162349 20051
rect 162259 19961 162287 19989
rect 162321 19961 162349 19989
rect 177619 20147 177647 20175
rect 177681 20147 177709 20175
rect 177619 20085 177647 20113
rect 177681 20085 177709 20113
rect 177619 20023 177647 20051
rect 177681 20023 177709 20051
rect 177619 19961 177647 19989
rect 177681 19961 177709 19989
rect 192979 20147 193007 20175
rect 193041 20147 193069 20175
rect 192979 20085 193007 20113
rect 193041 20085 193069 20113
rect 192979 20023 193007 20051
rect 193041 20023 193069 20051
rect 192979 19961 193007 19989
rect 193041 19961 193069 19989
rect 208339 20147 208367 20175
rect 208401 20147 208429 20175
rect 208339 20085 208367 20113
rect 208401 20085 208429 20113
rect 208339 20023 208367 20051
rect 208401 20023 208429 20051
rect 208339 19961 208367 19989
rect 208401 19961 208429 19989
rect 223699 20147 223727 20175
rect 223761 20147 223789 20175
rect 223699 20085 223727 20113
rect 223761 20085 223789 20113
rect 223699 20023 223727 20051
rect 223761 20023 223789 20051
rect 223699 19961 223727 19989
rect 223761 19961 223789 19989
rect 239059 20147 239087 20175
rect 239121 20147 239149 20175
rect 239059 20085 239087 20113
rect 239121 20085 239149 20113
rect 239059 20023 239087 20051
rect 239121 20023 239149 20051
rect 239059 19961 239087 19989
rect 239121 19961 239149 19989
rect 254419 20147 254447 20175
rect 254481 20147 254509 20175
rect 254419 20085 254447 20113
rect 254481 20085 254509 20113
rect 254419 20023 254447 20051
rect 254481 20023 254509 20051
rect 254419 19961 254447 19989
rect 254481 19961 254509 19989
rect 269779 20147 269807 20175
rect 269841 20147 269869 20175
rect 269779 20085 269807 20113
rect 269841 20085 269869 20113
rect 269779 20023 269807 20051
rect 269841 20023 269869 20051
rect 269779 19961 269807 19989
rect 269841 19961 269869 19989
rect 158217 14147 158245 14175
rect 158279 14147 158307 14175
rect 158341 14147 158369 14175
rect 158403 14147 158431 14175
rect 158217 14085 158245 14113
rect 158279 14085 158307 14113
rect 158341 14085 158369 14113
rect 158403 14085 158431 14113
rect 158217 14023 158245 14051
rect 158279 14023 158307 14051
rect 158341 14023 158369 14051
rect 158403 14023 158431 14051
rect 158217 13961 158245 13989
rect 158279 13961 158307 13989
rect 158341 13961 158369 13989
rect 158403 13961 158431 13989
rect 169939 14147 169967 14175
rect 170001 14147 170029 14175
rect 169939 14085 169967 14113
rect 170001 14085 170029 14113
rect 169939 14023 169967 14051
rect 170001 14023 170029 14051
rect 169939 13961 169967 13989
rect 170001 13961 170029 13989
rect 185299 14147 185327 14175
rect 185361 14147 185389 14175
rect 185299 14085 185327 14113
rect 185361 14085 185389 14113
rect 185299 14023 185327 14051
rect 185361 14023 185389 14051
rect 185299 13961 185327 13989
rect 185361 13961 185389 13989
rect 200659 14147 200687 14175
rect 200721 14147 200749 14175
rect 200659 14085 200687 14113
rect 200721 14085 200749 14113
rect 200659 14023 200687 14051
rect 200721 14023 200749 14051
rect 200659 13961 200687 13989
rect 200721 13961 200749 13989
rect 216019 14147 216047 14175
rect 216081 14147 216109 14175
rect 216019 14085 216047 14113
rect 216081 14085 216109 14113
rect 216019 14023 216047 14051
rect 216081 14023 216109 14051
rect 216019 13961 216047 13989
rect 216081 13961 216109 13989
rect 231379 14147 231407 14175
rect 231441 14147 231469 14175
rect 231379 14085 231407 14113
rect 231441 14085 231469 14113
rect 231379 14023 231407 14051
rect 231441 14023 231469 14051
rect 231379 13961 231407 13989
rect 231441 13961 231469 13989
rect 246739 14147 246767 14175
rect 246801 14147 246829 14175
rect 246739 14085 246767 14113
rect 246801 14085 246829 14113
rect 246739 14023 246767 14051
rect 246801 14023 246829 14051
rect 246739 13961 246767 13989
rect 246801 13961 246829 13989
rect 262099 14147 262127 14175
rect 262161 14147 262189 14175
rect 262099 14085 262127 14113
rect 262161 14085 262189 14113
rect 262099 14023 262127 14051
rect 262161 14023 262189 14051
rect 262099 13961 262127 13989
rect 262161 13961 262189 13989
rect 162259 11147 162287 11175
rect 162321 11147 162349 11175
rect 162259 11085 162287 11113
rect 162321 11085 162349 11113
rect 162259 11023 162287 11051
rect 162321 11023 162349 11051
rect 162259 10961 162287 10989
rect 162321 10961 162349 10989
rect 177619 11147 177647 11175
rect 177681 11147 177709 11175
rect 177619 11085 177647 11113
rect 177681 11085 177709 11113
rect 177619 11023 177647 11051
rect 177681 11023 177709 11051
rect 177619 10961 177647 10989
rect 177681 10961 177709 10989
rect 192979 11147 193007 11175
rect 193041 11147 193069 11175
rect 192979 11085 193007 11113
rect 193041 11085 193069 11113
rect 192979 11023 193007 11051
rect 193041 11023 193069 11051
rect 192979 10961 193007 10989
rect 193041 10961 193069 10989
rect 208339 11147 208367 11175
rect 208401 11147 208429 11175
rect 208339 11085 208367 11113
rect 208401 11085 208429 11113
rect 208339 11023 208367 11051
rect 208401 11023 208429 11051
rect 208339 10961 208367 10989
rect 208401 10961 208429 10989
rect 223699 11147 223727 11175
rect 223761 11147 223789 11175
rect 223699 11085 223727 11113
rect 223761 11085 223789 11113
rect 223699 11023 223727 11051
rect 223761 11023 223789 11051
rect 223699 10961 223727 10989
rect 223761 10961 223789 10989
rect 239059 11147 239087 11175
rect 239121 11147 239149 11175
rect 239059 11085 239087 11113
rect 239121 11085 239149 11113
rect 239059 11023 239087 11051
rect 239121 11023 239149 11051
rect 239059 10961 239087 10989
rect 239121 10961 239149 10989
rect 254419 11147 254447 11175
rect 254481 11147 254509 11175
rect 254419 11085 254447 11113
rect 254481 11085 254509 11113
rect 254419 11023 254447 11051
rect 254481 11023 254509 11051
rect 254419 10961 254447 10989
rect 254481 10961 254509 10989
rect 269779 11147 269807 11175
rect 269841 11147 269869 11175
rect 269779 11085 269807 11113
rect 269841 11085 269869 11113
rect 269779 11023 269807 11051
rect 269841 11023 269869 11051
rect 269779 10961 269807 10989
rect 269841 10961 269869 10989
rect 158217 5147 158245 5175
rect 158279 5147 158307 5175
rect 158341 5147 158369 5175
rect 158403 5147 158431 5175
rect 158217 5085 158245 5113
rect 158279 5085 158307 5113
rect 158341 5085 158369 5113
rect 158403 5085 158431 5113
rect 158217 5023 158245 5051
rect 158279 5023 158307 5051
rect 158341 5023 158369 5051
rect 158403 5023 158431 5051
rect 158217 4961 158245 4989
rect 158279 4961 158307 4989
rect 158341 4961 158369 4989
rect 158403 4961 158431 4989
rect 158217 -588 158245 -560
rect 158279 -588 158307 -560
rect 158341 -588 158369 -560
rect 158403 -588 158431 -560
rect 158217 -650 158245 -622
rect 158279 -650 158307 -622
rect 158341 -650 158369 -622
rect 158403 -650 158431 -622
rect 158217 -712 158245 -684
rect 158279 -712 158307 -684
rect 158341 -712 158369 -684
rect 158403 -712 158431 -684
rect 158217 -774 158245 -746
rect 158279 -774 158307 -746
rect 158341 -774 158369 -746
rect 158403 -774 158431 -746
rect 171717 2147 171745 2175
rect 171779 2147 171807 2175
rect 171841 2147 171869 2175
rect 171903 2147 171931 2175
rect 171717 2085 171745 2113
rect 171779 2085 171807 2113
rect 171841 2085 171869 2113
rect 171903 2085 171931 2113
rect 171717 2023 171745 2051
rect 171779 2023 171807 2051
rect 171841 2023 171869 2051
rect 171903 2023 171931 2051
rect 171717 1961 171745 1989
rect 171779 1961 171807 1989
rect 171841 1961 171869 1989
rect 171903 1961 171931 1989
rect 171717 -108 171745 -80
rect 171779 -108 171807 -80
rect 171841 -108 171869 -80
rect 171903 -108 171931 -80
rect 171717 -170 171745 -142
rect 171779 -170 171807 -142
rect 171841 -170 171869 -142
rect 171903 -170 171931 -142
rect 171717 -232 171745 -204
rect 171779 -232 171807 -204
rect 171841 -232 171869 -204
rect 171903 -232 171931 -204
rect 171717 -294 171745 -266
rect 171779 -294 171807 -266
rect 171841 -294 171869 -266
rect 171903 -294 171931 -266
rect 173577 5147 173605 5175
rect 173639 5147 173667 5175
rect 173701 5147 173729 5175
rect 173763 5147 173791 5175
rect 173577 5085 173605 5113
rect 173639 5085 173667 5113
rect 173701 5085 173729 5113
rect 173763 5085 173791 5113
rect 173577 5023 173605 5051
rect 173639 5023 173667 5051
rect 173701 5023 173729 5051
rect 173763 5023 173791 5051
rect 173577 4961 173605 4989
rect 173639 4961 173667 4989
rect 173701 4961 173729 4989
rect 173763 4961 173791 4989
rect 173577 -588 173605 -560
rect 173639 -588 173667 -560
rect 173701 -588 173729 -560
rect 173763 -588 173791 -560
rect 173577 -650 173605 -622
rect 173639 -650 173667 -622
rect 173701 -650 173729 -622
rect 173763 -650 173791 -622
rect 173577 -712 173605 -684
rect 173639 -712 173667 -684
rect 173701 -712 173729 -684
rect 173763 -712 173791 -684
rect 173577 -774 173605 -746
rect 173639 -774 173667 -746
rect 173701 -774 173729 -746
rect 173763 -774 173791 -746
rect 187077 2147 187105 2175
rect 187139 2147 187167 2175
rect 187201 2147 187229 2175
rect 187263 2147 187291 2175
rect 187077 2085 187105 2113
rect 187139 2085 187167 2113
rect 187201 2085 187229 2113
rect 187263 2085 187291 2113
rect 187077 2023 187105 2051
rect 187139 2023 187167 2051
rect 187201 2023 187229 2051
rect 187263 2023 187291 2051
rect 187077 1961 187105 1989
rect 187139 1961 187167 1989
rect 187201 1961 187229 1989
rect 187263 1961 187291 1989
rect 187077 -108 187105 -80
rect 187139 -108 187167 -80
rect 187201 -108 187229 -80
rect 187263 -108 187291 -80
rect 187077 -170 187105 -142
rect 187139 -170 187167 -142
rect 187201 -170 187229 -142
rect 187263 -170 187291 -142
rect 187077 -232 187105 -204
rect 187139 -232 187167 -204
rect 187201 -232 187229 -204
rect 187263 -232 187291 -204
rect 187077 -294 187105 -266
rect 187139 -294 187167 -266
rect 187201 -294 187229 -266
rect 187263 -294 187291 -266
rect 188937 5147 188965 5175
rect 188999 5147 189027 5175
rect 189061 5147 189089 5175
rect 189123 5147 189151 5175
rect 188937 5085 188965 5113
rect 188999 5085 189027 5113
rect 189061 5085 189089 5113
rect 189123 5085 189151 5113
rect 188937 5023 188965 5051
rect 188999 5023 189027 5051
rect 189061 5023 189089 5051
rect 189123 5023 189151 5051
rect 188937 4961 188965 4989
rect 188999 4961 189027 4989
rect 189061 4961 189089 4989
rect 189123 4961 189151 4989
rect 188937 -588 188965 -560
rect 188999 -588 189027 -560
rect 189061 -588 189089 -560
rect 189123 -588 189151 -560
rect 188937 -650 188965 -622
rect 188999 -650 189027 -622
rect 189061 -650 189089 -622
rect 189123 -650 189151 -622
rect 188937 -712 188965 -684
rect 188999 -712 189027 -684
rect 189061 -712 189089 -684
rect 189123 -712 189151 -684
rect 188937 -774 188965 -746
rect 188999 -774 189027 -746
rect 189061 -774 189089 -746
rect 189123 -774 189151 -746
rect 202437 2147 202465 2175
rect 202499 2147 202527 2175
rect 202561 2147 202589 2175
rect 202623 2147 202651 2175
rect 202437 2085 202465 2113
rect 202499 2085 202527 2113
rect 202561 2085 202589 2113
rect 202623 2085 202651 2113
rect 202437 2023 202465 2051
rect 202499 2023 202527 2051
rect 202561 2023 202589 2051
rect 202623 2023 202651 2051
rect 202437 1961 202465 1989
rect 202499 1961 202527 1989
rect 202561 1961 202589 1989
rect 202623 1961 202651 1989
rect 202437 -108 202465 -80
rect 202499 -108 202527 -80
rect 202561 -108 202589 -80
rect 202623 -108 202651 -80
rect 202437 -170 202465 -142
rect 202499 -170 202527 -142
rect 202561 -170 202589 -142
rect 202623 -170 202651 -142
rect 202437 -232 202465 -204
rect 202499 -232 202527 -204
rect 202561 -232 202589 -204
rect 202623 -232 202651 -204
rect 202437 -294 202465 -266
rect 202499 -294 202527 -266
rect 202561 -294 202589 -266
rect 202623 -294 202651 -266
rect 204297 5147 204325 5175
rect 204359 5147 204387 5175
rect 204421 5147 204449 5175
rect 204483 5147 204511 5175
rect 204297 5085 204325 5113
rect 204359 5085 204387 5113
rect 204421 5085 204449 5113
rect 204483 5085 204511 5113
rect 204297 5023 204325 5051
rect 204359 5023 204387 5051
rect 204421 5023 204449 5051
rect 204483 5023 204511 5051
rect 204297 4961 204325 4989
rect 204359 4961 204387 4989
rect 204421 4961 204449 4989
rect 204483 4961 204511 4989
rect 204297 -588 204325 -560
rect 204359 -588 204387 -560
rect 204421 -588 204449 -560
rect 204483 -588 204511 -560
rect 204297 -650 204325 -622
rect 204359 -650 204387 -622
rect 204421 -650 204449 -622
rect 204483 -650 204511 -622
rect 204297 -712 204325 -684
rect 204359 -712 204387 -684
rect 204421 -712 204449 -684
rect 204483 -712 204511 -684
rect 204297 -774 204325 -746
rect 204359 -774 204387 -746
rect 204421 -774 204449 -746
rect 204483 -774 204511 -746
rect 217797 2147 217825 2175
rect 217859 2147 217887 2175
rect 217921 2147 217949 2175
rect 217983 2147 218011 2175
rect 217797 2085 217825 2113
rect 217859 2085 217887 2113
rect 217921 2085 217949 2113
rect 217983 2085 218011 2113
rect 217797 2023 217825 2051
rect 217859 2023 217887 2051
rect 217921 2023 217949 2051
rect 217983 2023 218011 2051
rect 217797 1961 217825 1989
rect 217859 1961 217887 1989
rect 217921 1961 217949 1989
rect 217983 1961 218011 1989
rect 217797 -108 217825 -80
rect 217859 -108 217887 -80
rect 217921 -108 217949 -80
rect 217983 -108 218011 -80
rect 217797 -170 217825 -142
rect 217859 -170 217887 -142
rect 217921 -170 217949 -142
rect 217983 -170 218011 -142
rect 217797 -232 217825 -204
rect 217859 -232 217887 -204
rect 217921 -232 217949 -204
rect 217983 -232 218011 -204
rect 217797 -294 217825 -266
rect 217859 -294 217887 -266
rect 217921 -294 217949 -266
rect 217983 -294 218011 -266
rect 219657 5147 219685 5175
rect 219719 5147 219747 5175
rect 219781 5147 219809 5175
rect 219843 5147 219871 5175
rect 219657 5085 219685 5113
rect 219719 5085 219747 5113
rect 219781 5085 219809 5113
rect 219843 5085 219871 5113
rect 219657 5023 219685 5051
rect 219719 5023 219747 5051
rect 219781 5023 219809 5051
rect 219843 5023 219871 5051
rect 219657 4961 219685 4989
rect 219719 4961 219747 4989
rect 219781 4961 219809 4989
rect 219843 4961 219871 4989
rect 219657 -588 219685 -560
rect 219719 -588 219747 -560
rect 219781 -588 219809 -560
rect 219843 -588 219871 -560
rect 219657 -650 219685 -622
rect 219719 -650 219747 -622
rect 219781 -650 219809 -622
rect 219843 -650 219871 -622
rect 219657 -712 219685 -684
rect 219719 -712 219747 -684
rect 219781 -712 219809 -684
rect 219843 -712 219871 -684
rect 219657 -774 219685 -746
rect 219719 -774 219747 -746
rect 219781 -774 219809 -746
rect 219843 -774 219871 -746
rect 233157 2147 233185 2175
rect 233219 2147 233247 2175
rect 233281 2147 233309 2175
rect 233343 2147 233371 2175
rect 233157 2085 233185 2113
rect 233219 2085 233247 2113
rect 233281 2085 233309 2113
rect 233343 2085 233371 2113
rect 233157 2023 233185 2051
rect 233219 2023 233247 2051
rect 233281 2023 233309 2051
rect 233343 2023 233371 2051
rect 233157 1961 233185 1989
rect 233219 1961 233247 1989
rect 233281 1961 233309 1989
rect 233343 1961 233371 1989
rect 233157 -108 233185 -80
rect 233219 -108 233247 -80
rect 233281 -108 233309 -80
rect 233343 -108 233371 -80
rect 233157 -170 233185 -142
rect 233219 -170 233247 -142
rect 233281 -170 233309 -142
rect 233343 -170 233371 -142
rect 233157 -232 233185 -204
rect 233219 -232 233247 -204
rect 233281 -232 233309 -204
rect 233343 -232 233371 -204
rect 233157 -294 233185 -266
rect 233219 -294 233247 -266
rect 233281 -294 233309 -266
rect 233343 -294 233371 -266
rect 235017 5147 235045 5175
rect 235079 5147 235107 5175
rect 235141 5147 235169 5175
rect 235203 5147 235231 5175
rect 235017 5085 235045 5113
rect 235079 5085 235107 5113
rect 235141 5085 235169 5113
rect 235203 5085 235231 5113
rect 235017 5023 235045 5051
rect 235079 5023 235107 5051
rect 235141 5023 235169 5051
rect 235203 5023 235231 5051
rect 235017 4961 235045 4989
rect 235079 4961 235107 4989
rect 235141 4961 235169 4989
rect 235203 4961 235231 4989
rect 235017 -588 235045 -560
rect 235079 -588 235107 -560
rect 235141 -588 235169 -560
rect 235203 -588 235231 -560
rect 235017 -650 235045 -622
rect 235079 -650 235107 -622
rect 235141 -650 235169 -622
rect 235203 -650 235231 -622
rect 235017 -712 235045 -684
rect 235079 -712 235107 -684
rect 235141 -712 235169 -684
rect 235203 -712 235231 -684
rect 235017 -774 235045 -746
rect 235079 -774 235107 -746
rect 235141 -774 235169 -746
rect 235203 -774 235231 -746
rect 248517 2147 248545 2175
rect 248579 2147 248607 2175
rect 248641 2147 248669 2175
rect 248703 2147 248731 2175
rect 248517 2085 248545 2113
rect 248579 2085 248607 2113
rect 248641 2085 248669 2113
rect 248703 2085 248731 2113
rect 248517 2023 248545 2051
rect 248579 2023 248607 2051
rect 248641 2023 248669 2051
rect 248703 2023 248731 2051
rect 248517 1961 248545 1989
rect 248579 1961 248607 1989
rect 248641 1961 248669 1989
rect 248703 1961 248731 1989
rect 248517 -108 248545 -80
rect 248579 -108 248607 -80
rect 248641 -108 248669 -80
rect 248703 -108 248731 -80
rect 248517 -170 248545 -142
rect 248579 -170 248607 -142
rect 248641 -170 248669 -142
rect 248703 -170 248731 -142
rect 248517 -232 248545 -204
rect 248579 -232 248607 -204
rect 248641 -232 248669 -204
rect 248703 -232 248731 -204
rect 248517 -294 248545 -266
rect 248579 -294 248607 -266
rect 248641 -294 248669 -266
rect 248703 -294 248731 -266
rect 250377 5147 250405 5175
rect 250439 5147 250467 5175
rect 250501 5147 250529 5175
rect 250563 5147 250591 5175
rect 250377 5085 250405 5113
rect 250439 5085 250467 5113
rect 250501 5085 250529 5113
rect 250563 5085 250591 5113
rect 250377 5023 250405 5051
rect 250439 5023 250467 5051
rect 250501 5023 250529 5051
rect 250563 5023 250591 5051
rect 250377 4961 250405 4989
rect 250439 4961 250467 4989
rect 250501 4961 250529 4989
rect 250563 4961 250591 4989
rect 250377 -588 250405 -560
rect 250439 -588 250467 -560
rect 250501 -588 250529 -560
rect 250563 -588 250591 -560
rect 250377 -650 250405 -622
rect 250439 -650 250467 -622
rect 250501 -650 250529 -622
rect 250563 -650 250591 -622
rect 250377 -712 250405 -684
rect 250439 -712 250467 -684
rect 250501 -712 250529 -684
rect 250563 -712 250591 -684
rect 250377 -774 250405 -746
rect 250439 -774 250467 -746
rect 250501 -774 250529 -746
rect 250563 -774 250591 -746
rect 263877 2147 263905 2175
rect 263939 2147 263967 2175
rect 264001 2147 264029 2175
rect 264063 2147 264091 2175
rect 263877 2085 263905 2113
rect 263939 2085 263967 2113
rect 264001 2085 264029 2113
rect 264063 2085 264091 2113
rect 263877 2023 263905 2051
rect 263939 2023 263967 2051
rect 264001 2023 264029 2051
rect 264063 2023 264091 2051
rect 263877 1961 263905 1989
rect 263939 1961 263967 1989
rect 264001 1961 264029 1989
rect 264063 1961 264091 1989
rect 263877 -108 263905 -80
rect 263939 -108 263967 -80
rect 264001 -108 264029 -80
rect 264063 -108 264091 -80
rect 263877 -170 263905 -142
rect 263939 -170 263967 -142
rect 264001 -170 264029 -142
rect 264063 -170 264091 -142
rect 263877 -232 263905 -204
rect 263939 -232 263967 -204
rect 264001 -232 264029 -204
rect 264063 -232 264091 -204
rect 263877 -294 263905 -266
rect 263939 -294 263967 -266
rect 264001 -294 264029 -266
rect 264063 -294 264091 -266
rect 265737 5147 265765 5175
rect 265799 5147 265827 5175
rect 265861 5147 265889 5175
rect 265923 5147 265951 5175
rect 265737 5085 265765 5113
rect 265799 5085 265827 5113
rect 265861 5085 265889 5113
rect 265923 5085 265951 5113
rect 265737 5023 265765 5051
rect 265799 5023 265827 5051
rect 265861 5023 265889 5051
rect 265923 5023 265951 5051
rect 265737 4961 265765 4989
rect 265799 4961 265827 4989
rect 265861 4961 265889 4989
rect 265923 4961 265951 4989
rect 279237 146023 279265 146051
rect 279299 146023 279327 146051
rect 279361 146023 279389 146051
rect 279423 146023 279451 146051
rect 279237 145961 279265 145989
rect 279299 145961 279327 145989
rect 279361 145961 279389 145989
rect 279423 145961 279451 145989
rect 279237 137147 279265 137175
rect 279299 137147 279327 137175
rect 279361 137147 279389 137175
rect 279423 137147 279451 137175
rect 279237 137085 279265 137113
rect 279299 137085 279327 137113
rect 279361 137085 279389 137113
rect 279423 137085 279451 137113
rect 279237 137023 279265 137051
rect 279299 137023 279327 137051
rect 279361 137023 279389 137051
rect 279423 137023 279451 137051
rect 279237 136961 279265 136989
rect 279299 136961 279327 136989
rect 279361 136961 279389 136989
rect 279423 136961 279451 136989
rect 279237 128147 279265 128175
rect 279299 128147 279327 128175
rect 279361 128147 279389 128175
rect 279423 128147 279451 128175
rect 279237 128085 279265 128113
rect 279299 128085 279327 128113
rect 279361 128085 279389 128113
rect 279423 128085 279451 128113
rect 279237 128023 279265 128051
rect 279299 128023 279327 128051
rect 279361 128023 279389 128051
rect 279423 128023 279451 128051
rect 279237 127961 279265 127989
rect 279299 127961 279327 127989
rect 279361 127961 279389 127989
rect 279423 127961 279451 127989
rect 279237 119147 279265 119175
rect 279299 119147 279327 119175
rect 279361 119147 279389 119175
rect 279423 119147 279451 119175
rect 279237 119085 279265 119113
rect 279299 119085 279327 119113
rect 279361 119085 279389 119113
rect 279423 119085 279451 119113
rect 279237 119023 279265 119051
rect 279299 119023 279327 119051
rect 279361 119023 279389 119051
rect 279423 119023 279451 119051
rect 279237 118961 279265 118989
rect 279299 118961 279327 118989
rect 279361 118961 279389 118989
rect 279423 118961 279451 118989
rect 279237 110147 279265 110175
rect 279299 110147 279327 110175
rect 279361 110147 279389 110175
rect 279423 110147 279451 110175
rect 279237 110085 279265 110113
rect 279299 110085 279327 110113
rect 279361 110085 279389 110113
rect 279423 110085 279451 110113
rect 279237 110023 279265 110051
rect 279299 110023 279327 110051
rect 279361 110023 279389 110051
rect 279423 110023 279451 110051
rect 279237 109961 279265 109989
rect 279299 109961 279327 109989
rect 279361 109961 279389 109989
rect 279423 109961 279451 109989
rect 279237 101147 279265 101175
rect 279299 101147 279327 101175
rect 279361 101147 279389 101175
rect 279423 101147 279451 101175
rect 279237 101085 279265 101113
rect 279299 101085 279327 101113
rect 279361 101085 279389 101113
rect 279423 101085 279451 101113
rect 279237 101023 279265 101051
rect 279299 101023 279327 101051
rect 279361 101023 279389 101051
rect 279423 101023 279451 101051
rect 279237 100961 279265 100989
rect 279299 100961 279327 100989
rect 279361 100961 279389 100989
rect 279423 100961 279451 100989
rect 279237 92147 279265 92175
rect 279299 92147 279327 92175
rect 279361 92147 279389 92175
rect 279423 92147 279451 92175
rect 279237 92085 279265 92113
rect 279299 92085 279327 92113
rect 279361 92085 279389 92113
rect 279423 92085 279451 92113
rect 279237 92023 279265 92051
rect 279299 92023 279327 92051
rect 279361 92023 279389 92051
rect 279423 92023 279451 92051
rect 279237 91961 279265 91989
rect 279299 91961 279327 91989
rect 279361 91961 279389 91989
rect 279423 91961 279451 91989
rect 279237 83147 279265 83175
rect 279299 83147 279327 83175
rect 279361 83147 279389 83175
rect 279423 83147 279451 83175
rect 279237 83085 279265 83113
rect 279299 83085 279327 83113
rect 279361 83085 279389 83113
rect 279423 83085 279451 83113
rect 279237 83023 279265 83051
rect 279299 83023 279327 83051
rect 279361 83023 279389 83051
rect 279423 83023 279451 83051
rect 279237 82961 279265 82989
rect 279299 82961 279327 82989
rect 279361 82961 279389 82989
rect 279423 82961 279451 82989
rect 279237 74147 279265 74175
rect 279299 74147 279327 74175
rect 279361 74147 279389 74175
rect 279423 74147 279451 74175
rect 279237 74085 279265 74113
rect 279299 74085 279327 74113
rect 279361 74085 279389 74113
rect 279423 74085 279451 74113
rect 279237 74023 279265 74051
rect 279299 74023 279327 74051
rect 279361 74023 279389 74051
rect 279423 74023 279451 74051
rect 279237 73961 279265 73989
rect 279299 73961 279327 73989
rect 279361 73961 279389 73989
rect 279423 73961 279451 73989
rect 279237 65147 279265 65175
rect 279299 65147 279327 65175
rect 279361 65147 279389 65175
rect 279423 65147 279451 65175
rect 279237 65085 279265 65113
rect 279299 65085 279327 65113
rect 279361 65085 279389 65113
rect 279423 65085 279451 65113
rect 279237 65023 279265 65051
rect 279299 65023 279327 65051
rect 279361 65023 279389 65051
rect 279423 65023 279451 65051
rect 279237 64961 279265 64989
rect 279299 64961 279327 64989
rect 279361 64961 279389 64989
rect 279423 64961 279451 64989
rect 279237 56147 279265 56175
rect 279299 56147 279327 56175
rect 279361 56147 279389 56175
rect 279423 56147 279451 56175
rect 279237 56085 279265 56113
rect 279299 56085 279327 56113
rect 279361 56085 279389 56113
rect 279423 56085 279451 56113
rect 279237 56023 279265 56051
rect 279299 56023 279327 56051
rect 279361 56023 279389 56051
rect 279423 56023 279451 56051
rect 279237 55961 279265 55989
rect 279299 55961 279327 55989
rect 279361 55961 279389 55989
rect 279423 55961 279451 55989
rect 279237 47147 279265 47175
rect 279299 47147 279327 47175
rect 279361 47147 279389 47175
rect 279423 47147 279451 47175
rect 279237 47085 279265 47113
rect 279299 47085 279327 47113
rect 279361 47085 279389 47113
rect 279423 47085 279451 47113
rect 279237 47023 279265 47051
rect 279299 47023 279327 47051
rect 279361 47023 279389 47051
rect 279423 47023 279451 47051
rect 279237 46961 279265 46989
rect 279299 46961 279327 46989
rect 279361 46961 279389 46989
rect 279423 46961 279451 46989
rect 279237 38147 279265 38175
rect 279299 38147 279327 38175
rect 279361 38147 279389 38175
rect 279423 38147 279451 38175
rect 279237 38085 279265 38113
rect 279299 38085 279327 38113
rect 279361 38085 279389 38113
rect 279423 38085 279451 38113
rect 279237 38023 279265 38051
rect 279299 38023 279327 38051
rect 279361 38023 279389 38051
rect 279423 38023 279451 38051
rect 279237 37961 279265 37989
rect 279299 37961 279327 37989
rect 279361 37961 279389 37989
rect 279423 37961 279451 37989
rect 279237 29147 279265 29175
rect 279299 29147 279327 29175
rect 279361 29147 279389 29175
rect 279423 29147 279451 29175
rect 279237 29085 279265 29113
rect 279299 29085 279327 29113
rect 279361 29085 279389 29113
rect 279423 29085 279451 29113
rect 279237 29023 279265 29051
rect 279299 29023 279327 29051
rect 279361 29023 279389 29051
rect 279423 29023 279451 29051
rect 279237 28961 279265 28989
rect 279299 28961 279327 28989
rect 279361 28961 279389 28989
rect 279423 28961 279451 28989
rect 279237 20147 279265 20175
rect 279299 20147 279327 20175
rect 279361 20147 279389 20175
rect 279423 20147 279451 20175
rect 279237 20085 279265 20113
rect 279299 20085 279327 20113
rect 279361 20085 279389 20113
rect 279423 20085 279451 20113
rect 279237 20023 279265 20051
rect 279299 20023 279327 20051
rect 279361 20023 279389 20051
rect 279423 20023 279451 20051
rect 279237 19961 279265 19989
rect 279299 19961 279327 19989
rect 279361 19961 279389 19989
rect 279423 19961 279451 19989
rect 279237 11147 279265 11175
rect 279299 11147 279327 11175
rect 279361 11147 279389 11175
rect 279423 11147 279451 11175
rect 279237 11085 279265 11113
rect 279299 11085 279327 11113
rect 279361 11085 279389 11113
rect 279423 11085 279451 11113
rect 279237 11023 279265 11051
rect 279299 11023 279327 11051
rect 279361 11023 279389 11051
rect 279423 11023 279451 11051
rect 279237 10961 279265 10989
rect 279299 10961 279327 10989
rect 279361 10961 279389 10989
rect 279423 10961 279451 10989
rect 265737 -588 265765 -560
rect 265799 -588 265827 -560
rect 265861 -588 265889 -560
rect 265923 -588 265951 -560
rect 265737 -650 265765 -622
rect 265799 -650 265827 -622
rect 265861 -650 265889 -622
rect 265923 -650 265951 -622
rect 265737 -712 265765 -684
rect 265799 -712 265827 -684
rect 265861 -712 265889 -684
rect 265923 -712 265951 -684
rect 265737 -774 265765 -746
rect 265799 -774 265827 -746
rect 265861 -774 265889 -746
rect 265923 -774 265951 -746
rect 279237 2147 279265 2175
rect 279299 2147 279327 2175
rect 279361 2147 279389 2175
rect 279423 2147 279451 2175
rect 279237 2085 279265 2113
rect 279299 2085 279327 2113
rect 279361 2085 279389 2113
rect 279423 2085 279451 2113
rect 279237 2023 279265 2051
rect 279299 2023 279327 2051
rect 279361 2023 279389 2051
rect 279423 2023 279451 2051
rect 279237 1961 279265 1989
rect 279299 1961 279327 1989
rect 279361 1961 279389 1989
rect 279423 1961 279451 1989
rect 279237 -108 279265 -80
rect 279299 -108 279327 -80
rect 279361 -108 279389 -80
rect 279423 -108 279451 -80
rect 279237 -170 279265 -142
rect 279299 -170 279327 -142
rect 279361 -170 279389 -142
rect 279423 -170 279451 -142
rect 279237 -232 279265 -204
rect 279299 -232 279327 -204
rect 279361 -232 279389 -204
rect 279423 -232 279451 -204
rect 279237 -294 279265 -266
rect 279299 -294 279327 -266
rect 279361 -294 279389 -266
rect 279423 -294 279451 -266
rect 281097 299058 281125 299086
rect 281159 299058 281187 299086
rect 281221 299058 281249 299086
rect 281283 299058 281311 299086
rect 281097 298996 281125 299024
rect 281159 298996 281187 299024
rect 281221 298996 281249 299024
rect 281283 298996 281311 299024
rect 281097 298934 281125 298962
rect 281159 298934 281187 298962
rect 281221 298934 281249 298962
rect 281283 298934 281311 298962
rect 281097 298872 281125 298900
rect 281159 298872 281187 298900
rect 281221 298872 281249 298900
rect 281283 298872 281311 298900
rect 281097 293147 281125 293175
rect 281159 293147 281187 293175
rect 281221 293147 281249 293175
rect 281283 293147 281311 293175
rect 281097 293085 281125 293113
rect 281159 293085 281187 293113
rect 281221 293085 281249 293113
rect 281283 293085 281311 293113
rect 281097 293023 281125 293051
rect 281159 293023 281187 293051
rect 281221 293023 281249 293051
rect 281283 293023 281311 293051
rect 281097 292961 281125 292989
rect 281159 292961 281187 292989
rect 281221 292961 281249 292989
rect 281283 292961 281311 292989
rect 281097 284147 281125 284175
rect 281159 284147 281187 284175
rect 281221 284147 281249 284175
rect 281283 284147 281311 284175
rect 281097 284085 281125 284113
rect 281159 284085 281187 284113
rect 281221 284085 281249 284113
rect 281283 284085 281311 284113
rect 281097 284023 281125 284051
rect 281159 284023 281187 284051
rect 281221 284023 281249 284051
rect 281283 284023 281311 284051
rect 281097 283961 281125 283989
rect 281159 283961 281187 283989
rect 281221 283961 281249 283989
rect 281283 283961 281311 283989
rect 281097 275147 281125 275175
rect 281159 275147 281187 275175
rect 281221 275147 281249 275175
rect 281283 275147 281311 275175
rect 281097 275085 281125 275113
rect 281159 275085 281187 275113
rect 281221 275085 281249 275113
rect 281283 275085 281311 275113
rect 281097 275023 281125 275051
rect 281159 275023 281187 275051
rect 281221 275023 281249 275051
rect 281283 275023 281311 275051
rect 281097 274961 281125 274989
rect 281159 274961 281187 274989
rect 281221 274961 281249 274989
rect 281283 274961 281311 274989
rect 281097 266147 281125 266175
rect 281159 266147 281187 266175
rect 281221 266147 281249 266175
rect 281283 266147 281311 266175
rect 281097 266085 281125 266113
rect 281159 266085 281187 266113
rect 281221 266085 281249 266113
rect 281283 266085 281311 266113
rect 281097 266023 281125 266051
rect 281159 266023 281187 266051
rect 281221 266023 281249 266051
rect 281283 266023 281311 266051
rect 281097 265961 281125 265989
rect 281159 265961 281187 265989
rect 281221 265961 281249 265989
rect 281283 265961 281311 265989
rect 281097 257147 281125 257175
rect 281159 257147 281187 257175
rect 281221 257147 281249 257175
rect 281283 257147 281311 257175
rect 281097 257085 281125 257113
rect 281159 257085 281187 257113
rect 281221 257085 281249 257113
rect 281283 257085 281311 257113
rect 281097 257023 281125 257051
rect 281159 257023 281187 257051
rect 281221 257023 281249 257051
rect 281283 257023 281311 257051
rect 281097 256961 281125 256989
rect 281159 256961 281187 256989
rect 281221 256961 281249 256989
rect 281283 256961 281311 256989
rect 281097 248147 281125 248175
rect 281159 248147 281187 248175
rect 281221 248147 281249 248175
rect 281283 248147 281311 248175
rect 281097 248085 281125 248113
rect 281159 248085 281187 248113
rect 281221 248085 281249 248113
rect 281283 248085 281311 248113
rect 281097 248023 281125 248051
rect 281159 248023 281187 248051
rect 281221 248023 281249 248051
rect 281283 248023 281311 248051
rect 281097 247961 281125 247989
rect 281159 247961 281187 247989
rect 281221 247961 281249 247989
rect 281283 247961 281311 247989
rect 281097 239147 281125 239175
rect 281159 239147 281187 239175
rect 281221 239147 281249 239175
rect 281283 239147 281311 239175
rect 281097 239085 281125 239113
rect 281159 239085 281187 239113
rect 281221 239085 281249 239113
rect 281283 239085 281311 239113
rect 281097 239023 281125 239051
rect 281159 239023 281187 239051
rect 281221 239023 281249 239051
rect 281283 239023 281311 239051
rect 281097 238961 281125 238989
rect 281159 238961 281187 238989
rect 281221 238961 281249 238989
rect 281283 238961 281311 238989
rect 281097 230147 281125 230175
rect 281159 230147 281187 230175
rect 281221 230147 281249 230175
rect 281283 230147 281311 230175
rect 281097 230085 281125 230113
rect 281159 230085 281187 230113
rect 281221 230085 281249 230113
rect 281283 230085 281311 230113
rect 281097 230023 281125 230051
rect 281159 230023 281187 230051
rect 281221 230023 281249 230051
rect 281283 230023 281311 230051
rect 281097 229961 281125 229989
rect 281159 229961 281187 229989
rect 281221 229961 281249 229989
rect 281283 229961 281311 229989
rect 281097 221147 281125 221175
rect 281159 221147 281187 221175
rect 281221 221147 281249 221175
rect 281283 221147 281311 221175
rect 281097 221085 281125 221113
rect 281159 221085 281187 221113
rect 281221 221085 281249 221113
rect 281283 221085 281311 221113
rect 281097 221023 281125 221051
rect 281159 221023 281187 221051
rect 281221 221023 281249 221051
rect 281283 221023 281311 221051
rect 281097 220961 281125 220989
rect 281159 220961 281187 220989
rect 281221 220961 281249 220989
rect 281283 220961 281311 220989
rect 281097 212147 281125 212175
rect 281159 212147 281187 212175
rect 281221 212147 281249 212175
rect 281283 212147 281311 212175
rect 281097 212085 281125 212113
rect 281159 212085 281187 212113
rect 281221 212085 281249 212113
rect 281283 212085 281311 212113
rect 281097 212023 281125 212051
rect 281159 212023 281187 212051
rect 281221 212023 281249 212051
rect 281283 212023 281311 212051
rect 281097 211961 281125 211989
rect 281159 211961 281187 211989
rect 281221 211961 281249 211989
rect 281283 211961 281311 211989
rect 281097 203147 281125 203175
rect 281159 203147 281187 203175
rect 281221 203147 281249 203175
rect 281283 203147 281311 203175
rect 281097 203085 281125 203113
rect 281159 203085 281187 203113
rect 281221 203085 281249 203113
rect 281283 203085 281311 203113
rect 281097 203023 281125 203051
rect 281159 203023 281187 203051
rect 281221 203023 281249 203051
rect 281283 203023 281311 203051
rect 281097 202961 281125 202989
rect 281159 202961 281187 202989
rect 281221 202961 281249 202989
rect 281283 202961 281311 202989
rect 281097 194147 281125 194175
rect 281159 194147 281187 194175
rect 281221 194147 281249 194175
rect 281283 194147 281311 194175
rect 281097 194085 281125 194113
rect 281159 194085 281187 194113
rect 281221 194085 281249 194113
rect 281283 194085 281311 194113
rect 281097 194023 281125 194051
rect 281159 194023 281187 194051
rect 281221 194023 281249 194051
rect 281283 194023 281311 194051
rect 281097 193961 281125 193989
rect 281159 193961 281187 193989
rect 281221 193961 281249 193989
rect 281283 193961 281311 193989
rect 281097 185147 281125 185175
rect 281159 185147 281187 185175
rect 281221 185147 281249 185175
rect 281283 185147 281311 185175
rect 281097 185085 281125 185113
rect 281159 185085 281187 185113
rect 281221 185085 281249 185113
rect 281283 185085 281311 185113
rect 281097 185023 281125 185051
rect 281159 185023 281187 185051
rect 281221 185023 281249 185051
rect 281283 185023 281311 185051
rect 281097 184961 281125 184989
rect 281159 184961 281187 184989
rect 281221 184961 281249 184989
rect 281283 184961 281311 184989
rect 281097 176147 281125 176175
rect 281159 176147 281187 176175
rect 281221 176147 281249 176175
rect 281283 176147 281311 176175
rect 281097 176085 281125 176113
rect 281159 176085 281187 176113
rect 281221 176085 281249 176113
rect 281283 176085 281311 176113
rect 281097 176023 281125 176051
rect 281159 176023 281187 176051
rect 281221 176023 281249 176051
rect 281283 176023 281311 176051
rect 281097 175961 281125 175989
rect 281159 175961 281187 175989
rect 281221 175961 281249 175989
rect 281283 175961 281311 175989
rect 281097 167147 281125 167175
rect 281159 167147 281187 167175
rect 281221 167147 281249 167175
rect 281283 167147 281311 167175
rect 281097 167085 281125 167113
rect 281159 167085 281187 167113
rect 281221 167085 281249 167113
rect 281283 167085 281311 167113
rect 281097 167023 281125 167051
rect 281159 167023 281187 167051
rect 281221 167023 281249 167051
rect 281283 167023 281311 167051
rect 281097 166961 281125 166989
rect 281159 166961 281187 166989
rect 281221 166961 281249 166989
rect 281283 166961 281311 166989
rect 281097 158147 281125 158175
rect 281159 158147 281187 158175
rect 281221 158147 281249 158175
rect 281283 158147 281311 158175
rect 281097 158085 281125 158113
rect 281159 158085 281187 158113
rect 281221 158085 281249 158113
rect 281283 158085 281311 158113
rect 281097 158023 281125 158051
rect 281159 158023 281187 158051
rect 281221 158023 281249 158051
rect 281283 158023 281311 158051
rect 281097 157961 281125 157989
rect 281159 157961 281187 157989
rect 281221 157961 281249 157989
rect 281283 157961 281311 157989
rect 281097 149147 281125 149175
rect 281159 149147 281187 149175
rect 281221 149147 281249 149175
rect 281283 149147 281311 149175
rect 281097 149085 281125 149113
rect 281159 149085 281187 149113
rect 281221 149085 281249 149113
rect 281283 149085 281311 149113
rect 281097 149023 281125 149051
rect 281159 149023 281187 149051
rect 281221 149023 281249 149051
rect 281283 149023 281311 149051
rect 281097 148961 281125 148989
rect 281159 148961 281187 148989
rect 281221 148961 281249 148989
rect 281283 148961 281311 148989
rect 281097 140147 281125 140175
rect 281159 140147 281187 140175
rect 281221 140147 281249 140175
rect 281283 140147 281311 140175
rect 281097 140085 281125 140113
rect 281159 140085 281187 140113
rect 281221 140085 281249 140113
rect 281283 140085 281311 140113
rect 281097 140023 281125 140051
rect 281159 140023 281187 140051
rect 281221 140023 281249 140051
rect 281283 140023 281311 140051
rect 281097 139961 281125 139989
rect 281159 139961 281187 139989
rect 281221 139961 281249 139989
rect 281283 139961 281311 139989
rect 281097 131147 281125 131175
rect 281159 131147 281187 131175
rect 281221 131147 281249 131175
rect 281283 131147 281311 131175
rect 281097 131085 281125 131113
rect 281159 131085 281187 131113
rect 281221 131085 281249 131113
rect 281283 131085 281311 131113
rect 281097 131023 281125 131051
rect 281159 131023 281187 131051
rect 281221 131023 281249 131051
rect 281283 131023 281311 131051
rect 281097 130961 281125 130989
rect 281159 130961 281187 130989
rect 281221 130961 281249 130989
rect 281283 130961 281311 130989
rect 281097 122147 281125 122175
rect 281159 122147 281187 122175
rect 281221 122147 281249 122175
rect 281283 122147 281311 122175
rect 281097 122085 281125 122113
rect 281159 122085 281187 122113
rect 281221 122085 281249 122113
rect 281283 122085 281311 122113
rect 281097 122023 281125 122051
rect 281159 122023 281187 122051
rect 281221 122023 281249 122051
rect 281283 122023 281311 122051
rect 281097 121961 281125 121989
rect 281159 121961 281187 121989
rect 281221 121961 281249 121989
rect 281283 121961 281311 121989
rect 281097 113147 281125 113175
rect 281159 113147 281187 113175
rect 281221 113147 281249 113175
rect 281283 113147 281311 113175
rect 281097 113085 281125 113113
rect 281159 113085 281187 113113
rect 281221 113085 281249 113113
rect 281283 113085 281311 113113
rect 281097 113023 281125 113051
rect 281159 113023 281187 113051
rect 281221 113023 281249 113051
rect 281283 113023 281311 113051
rect 281097 112961 281125 112989
rect 281159 112961 281187 112989
rect 281221 112961 281249 112989
rect 281283 112961 281311 112989
rect 281097 104147 281125 104175
rect 281159 104147 281187 104175
rect 281221 104147 281249 104175
rect 281283 104147 281311 104175
rect 281097 104085 281125 104113
rect 281159 104085 281187 104113
rect 281221 104085 281249 104113
rect 281283 104085 281311 104113
rect 281097 104023 281125 104051
rect 281159 104023 281187 104051
rect 281221 104023 281249 104051
rect 281283 104023 281311 104051
rect 281097 103961 281125 103989
rect 281159 103961 281187 103989
rect 281221 103961 281249 103989
rect 281283 103961 281311 103989
rect 281097 95147 281125 95175
rect 281159 95147 281187 95175
rect 281221 95147 281249 95175
rect 281283 95147 281311 95175
rect 281097 95085 281125 95113
rect 281159 95085 281187 95113
rect 281221 95085 281249 95113
rect 281283 95085 281311 95113
rect 281097 95023 281125 95051
rect 281159 95023 281187 95051
rect 281221 95023 281249 95051
rect 281283 95023 281311 95051
rect 281097 94961 281125 94989
rect 281159 94961 281187 94989
rect 281221 94961 281249 94989
rect 281283 94961 281311 94989
rect 281097 86147 281125 86175
rect 281159 86147 281187 86175
rect 281221 86147 281249 86175
rect 281283 86147 281311 86175
rect 281097 86085 281125 86113
rect 281159 86085 281187 86113
rect 281221 86085 281249 86113
rect 281283 86085 281311 86113
rect 281097 86023 281125 86051
rect 281159 86023 281187 86051
rect 281221 86023 281249 86051
rect 281283 86023 281311 86051
rect 281097 85961 281125 85989
rect 281159 85961 281187 85989
rect 281221 85961 281249 85989
rect 281283 85961 281311 85989
rect 281097 77147 281125 77175
rect 281159 77147 281187 77175
rect 281221 77147 281249 77175
rect 281283 77147 281311 77175
rect 281097 77085 281125 77113
rect 281159 77085 281187 77113
rect 281221 77085 281249 77113
rect 281283 77085 281311 77113
rect 281097 77023 281125 77051
rect 281159 77023 281187 77051
rect 281221 77023 281249 77051
rect 281283 77023 281311 77051
rect 281097 76961 281125 76989
rect 281159 76961 281187 76989
rect 281221 76961 281249 76989
rect 281283 76961 281311 76989
rect 281097 68147 281125 68175
rect 281159 68147 281187 68175
rect 281221 68147 281249 68175
rect 281283 68147 281311 68175
rect 281097 68085 281125 68113
rect 281159 68085 281187 68113
rect 281221 68085 281249 68113
rect 281283 68085 281311 68113
rect 281097 68023 281125 68051
rect 281159 68023 281187 68051
rect 281221 68023 281249 68051
rect 281283 68023 281311 68051
rect 281097 67961 281125 67989
rect 281159 67961 281187 67989
rect 281221 67961 281249 67989
rect 281283 67961 281311 67989
rect 281097 59147 281125 59175
rect 281159 59147 281187 59175
rect 281221 59147 281249 59175
rect 281283 59147 281311 59175
rect 281097 59085 281125 59113
rect 281159 59085 281187 59113
rect 281221 59085 281249 59113
rect 281283 59085 281311 59113
rect 281097 59023 281125 59051
rect 281159 59023 281187 59051
rect 281221 59023 281249 59051
rect 281283 59023 281311 59051
rect 281097 58961 281125 58989
rect 281159 58961 281187 58989
rect 281221 58961 281249 58989
rect 281283 58961 281311 58989
rect 281097 50147 281125 50175
rect 281159 50147 281187 50175
rect 281221 50147 281249 50175
rect 281283 50147 281311 50175
rect 281097 50085 281125 50113
rect 281159 50085 281187 50113
rect 281221 50085 281249 50113
rect 281283 50085 281311 50113
rect 281097 50023 281125 50051
rect 281159 50023 281187 50051
rect 281221 50023 281249 50051
rect 281283 50023 281311 50051
rect 281097 49961 281125 49989
rect 281159 49961 281187 49989
rect 281221 49961 281249 49989
rect 281283 49961 281311 49989
rect 281097 41147 281125 41175
rect 281159 41147 281187 41175
rect 281221 41147 281249 41175
rect 281283 41147 281311 41175
rect 281097 41085 281125 41113
rect 281159 41085 281187 41113
rect 281221 41085 281249 41113
rect 281283 41085 281311 41113
rect 281097 41023 281125 41051
rect 281159 41023 281187 41051
rect 281221 41023 281249 41051
rect 281283 41023 281311 41051
rect 281097 40961 281125 40989
rect 281159 40961 281187 40989
rect 281221 40961 281249 40989
rect 281283 40961 281311 40989
rect 281097 32147 281125 32175
rect 281159 32147 281187 32175
rect 281221 32147 281249 32175
rect 281283 32147 281311 32175
rect 281097 32085 281125 32113
rect 281159 32085 281187 32113
rect 281221 32085 281249 32113
rect 281283 32085 281311 32113
rect 281097 32023 281125 32051
rect 281159 32023 281187 32051
rect 281221 32023 281249 32051
rect 281283 32023 281311 32051
rect 281097 31961 281125 31989
rect 281159 31961 281187 31989
rect 281221 31961 281249 31989
rect 281283 31961 281311 31989
rect 281097 23147 281125 23175
rect 281159 23147 281187 23175
rect 281221 23147 281249 23175
rect 281283 23147 281311 23175
rect 281097 23085 281125 23113
rect 281159 23085 281187 23113
rect 281221 23085 281249 23113
rect 281283 23085 281311 23113
rect 281097 23023 281125 23051
rect 281159 23023 281187 23051
rect 281221 23023 281249 23051
rect 281283 23023 281311 23051
rect 281097 22961 281125 22989
rect 281159 22961 281187 22989
rect 281221 22961 281249 22989
rect 281283 22961 281311 22989
rect 281097 14147 281125 14175
rect 281159 14147 281187 14175
rect 281221 14147 281249 14175
rect 281283 14147 281311 14175
rect 281097 14085 281125 14113
rect 281159 14085 281187 14113
rect 281221 14085 281249 14113
rect 281283 14085 281311 14113
rect 281097 14023 281125 14051
rect 281159 14023 281187 14051
rect 281221 14023 281249 14051
rect 281283 14023 281311 14051
rect 281097 13961 281125 13989
rect 281159 13961 281187 13989
rect 281221 13961 281249 13989
rect 281283 13961 281311 13989
rect 281097 5147 281125 5175
rect 281159 5147 281187 5175
rect 281221 5147 281249 5175
rect 281283 5147 281311 5175
rect 281097 5085 281125 5113
rect 281159 5085 281187 5113
rect 281221 5085 281249 5113
rect 281283 5085 281311 5113
rect 281097 5023 281125 5051
rect 281159 5023 281187 5051
rect 281221 5023 281249 5051
rect 281283 5023 281311 5051
rect 281097 4961 281125 4989
rect 281159 4961 281187 4989
rect 281221 4961 281249 4989
rect 281283 4961 281311 4989
rect 281097 -588 281125 -560
rect 281159 -588 281187 -560
rect 281221 -588 281249 -560
rect 281283 -588 281311 -560
rect 281097 -650 281125 -622
rect 281159 -650 281187 -622
rect 281221 -650 281249 -622
rect 281283 -650 281311 -622
rect 281097 -712 281125 -684
rect 281159 -712 281187 -684
rect 281221 -712 281249 -684
rect 281283 -712 281311 -684
rect 281097 -774 281125 -746
rect 281159 -774 281187 -746
rect 281221 -774 281249 -746
rect 281283 -774 281311 -746
rect 294597 298578 294625 298606
rect 294659 298578 294687 298606
rect 294721 298578 294749 298606
rect 294783 298578 294811 298606
rect 294597 298516 294625 298544
rect 294659 298516 294687 298544
rect 294721 298516 294749 298544
rect 294783 298516 294811 298544
rect 294597 298454 294625 298482
rect 294659 298454 294687 298482
rect 294721 298454 294749 298482
rect 294783 298454 294811 298482
rect 294597 298392 294625 298420
rect 294659 298392 294687 298420
rect 294721 298392 294749 298420
rect 294783 298392 294811 298420
rect 294597 290147 294625 290175
rect 294659 290147 294687 290175
rect 294721 290147 294749 290175
rect 294783 290147 294811 290175
rect 294597 290085 294625 290113
rect 294659 290085 294687 290113
rect 294721 290085 294749 290113
rect 294783 290085 294811 290113
rect 294597 290023 294625 290051
rect 294659 290023 294687 290051
rect 294721 290023 294749 290051
rect 294783 290023 294811 290051
rect 294597 289961 294625 289989
rect 294659 289961 294687 289989
rect 294721 289961 294749 289989
rect 294783 289961 294811 289989
rect 294597 281147 294625 281175
rect 294659 281147 294687 281175
rect 294721 281147 294749 281175
rect 294783 281147 294811 281175
rect 294597 281085 294625 281113
rect 294659 281085 294687 281113
rect 294721 281085 294749 281113
rect 294783 281085 294811 281113
rect 296457 299058 296485 299086
rect 296519 299058 296547 299086
rect 296581 299058 296609 299086
rect 296643 299058 296671 299086
rect 296457 298996 296485 299024
rect 296519 298996 296547 299024
rect 296581 298996 296609 299024
rect 296643 298996 296671 299024
rect 296457 298934 296485 298962
rect 296519 298934 296547 298962
rect 296581 298934 296609 298962
rect 296643 298934 296671 298962
rect 296457 298872 296485 298900
rect 296519 298872 296547 298900
rect 296581 298872 296609 298900
rect 296643 298872 296671 298900
rect 298728 299058 298756 299086
rect 298790 299058 298818 299086
rect 298852 299058 298880 299086
rect 298914 299058 298942 299086
rect 298728 298996 298756 299024
rect 298790 298996 298818 299024
rect 298852 298996 298880 299024
rect 298914 298996 298942 299024
rect 298728 298934 298756 298962
rect 298790 298934 298818 298962
rect 298852 298934 298880 298962
rect 298914 298934 298942 298962
rect 298728 298872 298756 298900
rect 298790 298872 298818 298900
rect 298852 298872 298880 298900
rect 298914 298872 298942 298900
rect 296457 293147 296485 293175
rect 296519 293147 296547 293175
rect 296581 293147 296609 293175
rect 296643 293147 296671 293175
rect 296457 293085 296485 293113
rect 296519 293085 296547 293113
rect 296581 293085 296609 293113
rect 296643 293085 296671 293113
rect 296457 293023 296485 293051
rect 296519 293023 296547 293051
rect 296581 293023 296609 293051
rect 296643 293023 296671 293051
rect 296457 292961 296485 292989
rect 296519 292961 296547 292989
rect 296581 292961 296609 292989
rect 296643 292961 296671 292989
rect 296457 284147 296485 284175
rect 296519 284147 296547 284175
rect 296581 284147 296609 284175
rect 296643 284147 296671 284175
rect 296457 284085 296485 284113
rect 296519 284085 296547 284113
rect 296581 284085 296609 284113
rect 296643 284085 296671 284113
rect 296457 284023 296485 284051
rect 296519 284023 296547 284051
rect 296581 284023 296609 284051
rect 296643 284023 296671 284051
rect 296457 283961 296485 283989
rect 296519 283961 296547 283989
rect 296581 283961 296609 283989
rect 296643 283961 296671 283989
rect 294597 281023 294625 281051
rect 294659 281023 294687 281051
rect 294721 281023 294749 281051
rect 294783 281023 294811 281051
rect 294597 280961 294625 280989
rect 294659 280961 294687 280989
rect 294721 280961 294749 280989
rect 294783 280961 294811 280989
rect 294597 272147 294625 272175
rect 294659 272147 294687 272175
rect 294721 272147 294749 272175
rect 294783 272147 294811 272175
rect 294597 272085 294625 272113
rect 294659 272085 294687 272113
rect 294721 272085 294749 272113
rect 294783 272085 294811 272113
rect 294597 272023 294625 272051
rect 294659 272023 294687 272051
rect 294721 272023 294749 272051
rect 294783 272023 294811 272051
rect 294597 271961 294625 271989
rect 294659 271961 294687 271989
rect 294721 271961 294749 271989
rect 294783 271961 294811 271989
rect 294597 263147 294625 263175
rect 294659 263147 294687 263175
rect 294721 263147 294749 263175
rect 294783 263147 294811 263175
rect 294597 263085 294625 263113
rect 294659 263085 294687 263113
rect 294721 263085 294749 263113
rect 294783 263085 294811 263113
rect 294597 263023 294625 263051
rect 294659 263023 294687 263051
rect 294721 263023 294749 263051
rect 294783 263023 294811 263051
rect 294597 262961 294625 262989
rect 294659 262961 294687 262989
rect 294721 262961 294749 262989
rect 294783 262961 294811 262989
rect 294597 254147 294625 254175
rect 294659 254147 294687 254175
rect 294721 254147 294749 254175
rect 294783 254147 294811 254175
rect 294597 254085 294625 254113
rect 294659 254085 294687 254113
rect 294721 254085 294749 254113
rect 294783 254085 294811 254113
rect 294597 254023 294625 254051
rect 294659 254023 294687 254051
rect 294721 254023 294749 254051
rect 294783 254023 294811 254051
rect 294597 253961 294625 253989
rect 294659 253961 294687 253989
rect 294721 253961 294749 253989
rect 294783 253961 294811 253989
rect 294597 245147 294625 245175
rect 294659 245147 294687 245175
rect 294721 245147 294749 245175
rect 294783 245147 294811 245175
rect 294597 245085 294625 245113
rect 294659 245085 294687 245113
rect 294721 245085 294749 245113
rect 294783 245085 294811 245113
rect 294597 245023 294625 245051
rect 294659 245023 294687 245051
rect 294721 245023 294749 245051
rect 294783 245023 294811 245051
rect 294597 244961 294625 244989
rect 294659 244961 294687 244989
rect 294721 244961 294749 244989
rect 294783 244961 294811 244989
rect 294597 236147 294625 236175
rect 294659 236147 294687 236175
rect 294721 236147 294749 236175
rect 294783 236147 294811 236175
rect 294597 236085 294625 236113
rect 294659 236085 294687 236113
rect 294721 236085 294749 236113
rect 294783 236085 294811 236113
rect 294597 236023 294625 236051
rect 294659 236023 294687 236051
rect 294721 236023 294749 236051
rect 294783 236023 294811 236051
rect 294597 235961 294625 235989
rect 294659 235961 294687 235989
rect 294721 235961 294749 235989
rect 294783 235961 294811 235989
rect 294597 227147 294625 227175
rect 294659 227147 294687 227175
rect 294721 227147 294749 227175
rect 294783 227147 294811 227175
rect 294597 227085 294625 227113
rect 294659 227085 294687 227113
rect 294721 227085 294749 227113
rect 294783 227085 294811 227113
rect 294597 227023 294625 227051
rect 294659 227023 294687 227051
rect 294721 227023 294749 227051
rect 294783 227023 294811 227051
rect 294597 226961 294625 226989
rect 294659 226961 294687 226989
rect 294721 226961 294749 226989
rect 294783 226961 294811 226989
rect 294597 218147 294625 218175
rect 294659 218147 294687 218175
rect 294721 218147 294749 218175
rect 294783 218147 294811 218175
rect 294597 218085 294625 218113
rect 294659 218085 294687 218113
rect 294721 218085 294749 218113
rect 294783 218085 294811 218113
rect 294597 218023 294625 218051
rect 294659 218023 294687 218051
rect 294721 218023 294749 218051
rect 294783 218023 294811 218051
rect 294597 217961 294625 217989
rect 294659 217961 294687 217989
rect 294721 217961 294749 217989
rect 294783 217961 294811 217989
rect 294597 209147 294625 209175
rect 294659 209147 294687 209175
rect 294721 209147 294749 209175
rect 294783 209147 294811 209175
rect 294597 209085 294625 209113
rect 294659 209085 294687 209113
rect 294721 209085 294749 209113
rect 294783 209085 294811 209113
rect 294597 209023 294625 209051
rect 294659 209023 294687 209051
rect 294721 209023 294749 209051
rect 294783 209023 294811 209051
rect 294597 208961 294625 208989
rect 294659 208961 294687 208989
rect 294721 208961 294749 208989
rect 294783 208961 294811 208989
rect 294597 200147 294625 200175
rect 294659 200147 294687 200175
rect 294721 200147 294749 200175
rect 294783 200147 294811 200175
rect 294597 200085 294625 200113
rect 294659 200085 294687 200113
rect 294721 200085 294749 200113
rect 294783 200085 294811 200113
rect 294597 200023 294625 200051
rect 294659 200023 294687 200051
rect 294721 200023 294749 200051
rect 294783 200023 294811 200051
rect 294597 199961 294625 199989
rect 294659 199961 294687 199989
rect 294721 199961 294749 199989
rect 294783 199961 294811 199989
rect 294597 191147 294625 191175
rect 294659 191147 294687 191175
rect 294721 191147 294749 191175
rect 294783 191147 294811 191175
rect 294597 191085 294625 191113
rect 294659 191085 294687 191113
rect 294721 191085 294749 191113
rect 294783 191085 294811 191113
rect 294597 191023 294625 191051
rect 294659 191023 294687 191051
rect 294721 191023 294749 191051
rect 294783 191023 294811 191051
rect 294597 190961 294625 190989
rect 294659 190961 294687 190989
rect 294721 190961 294749 190989
rect 294783 190961 294811 190989
rect 294597 182147 294625 182175
rect 294659 182147 294687 182175
rect 294721 182147 294749 182175
rect 294783 182147 294811 182175
rect 294597 182085 294625 182113
rect 294659 182085 294687 182113
rect 294721 182085 294749 182113
rect 294783 182085 294811 182113
rect 294597 182023 294625 182051
rect 294659 182023 294687 182051
rect 294721 182023 294749 182051
rect 294783 182023 294811 182051
rect 294597 181961 294625 181989
rect 294659 181961 294687 181989
rect 294721 181961 294749 181989
rect 294783 181961 294811 181989
rect 294597 173147 294625 173175
rect 294659 173147 294687 173175
rect 294721 173147 294749 173175
rect 294783 173147 294811 173175
rect 294597 173085 294625 173113
rect 294659 173085 294687 173113
rect 294721 173085 294749 173113
rect 294783 173085 294811 173113
rect 294597 173023 294625 173051
rect 294659 173023 294687 173051
rect 294721 173023 294749 173051
rect 294783 173023 294811 173051
rect 294597 172961 294625 172989
rect 294659 172961 294687 172989
rect 294721 172961 294749 172989
rect 294783 172961 294811 172989
rect 294597 164147 294625 164175
rect 294659 164147 294687 164175
rect 294721 164147 294749 164175
rect 294783 164147 294811 164175
rect 294597 164085 294625 164113
rect 294659 164085 294687 164113
rect 294721 164085 294749 164113
rect 294783 164085 294811 164113
rect 294597 164023 294625 164051
rect 294659 164023 294687 164051
rect 294721 164023 294749 164051
rect 294783 164023 294811 164051
rect 294597 163961 294625 163989
rect 294659 163961 294687 163989
rect 294721 163961 294749 163989
rect 294783 163961 294811 163989
rect 296457 275147 296485 275175
rect 296519 275147 296547 275175
rect 296581 275147 296609 275175
rect 296643 275147 296671 275175
rect 296457 275085 296485 275113
rect 296519 275085 296547 275113
rect 296581 275085 296609 275113
rect 296643 275085 296671 275113
rect 296457 275023 296485 275051
rect 296519 275023 296547 275051
rect 296581 275023 296609 275051
rect 296643 275023 296671 275051
rect 296457 274961 296485 274989
rect 296519 274961 296547 274989
rect 296581 274961 296609 274989
rect 296643 274961 296671 274989
rect 296457 266147 296485 266175
rect 296519 266147 296547 266175
rect 296581 266147 296609 266175
rect 296643 266147 296671 266175
rect 296457 266085 296485 266113
rect 296519 266085 296547 266113
rect 296581 266085 296609 266113
rect 296643 266085 296671 266113
rect 296457 266023 296485 266051
rect 296519 266023 296547 266051
rect 296581 266023 296609 266051
rect 296643 266023 296671 266051
rect 296457 265961 296485 265989
rect 296519 265961 296547 265989
rect 296581 265961 296609 265989
rect 296643 265961 296671 265989
rect 296457 257147 296485 257175
rect 296519 257147 296547 257175
rect 296581 257147 296609 257175
rect 296643 257147 296671 257175
rect 296457 257085 296485 257113
rect 296519 257085 296547 257113
rect 296581 257085 296609 257113
rect 296643 257085 296671 257113
rect 296457 257023 296485 257051
rect 296519 257023 296547 257051
rect 296581 257023 296609 257051
rect 296643 257023 296671 257051
rect 296457 256961 296485 256989
rect 296519 256961 296547 256989
rect 296581 256961 296609 256989
rect 296643 256961 296671 256989
rect 296457 248147 296485 248175
rect 296519 248147 296547 248175
rect 296581 248147 296609 248175
rect 296643 248147 296671 248175
rect 296457 248085 296485 248113
rect 296519 248085 296547 248113
rect 296581 248085 296609 248113
rect 296643 248085 296671 248113
rect 296457 248023 296485 248051
rect 296519 248023 296547 248051
rect 296581 248023 296609 248051
rect 296643 248023 296671 248051
rect 296457 247961 296485 247989
rect 296519 247961 296547 247989
rect 296581 247961 296609 247989
rect 296643 247961 296671 247989
rect 294597 155147 294625 155175
rect 294659 155147 294687 155175
rect 294721 155147 294749 155175
rect 294783 155147 294811 155175
rect 294597 155085 294625 155113
rect 294659 155085 294687 155113
rect 294721 155085 294749 155113
rect 294783 155085 294811 155113
rect 294597 155023 294625 155051
rect 294659 155023 294687 155051
rect 294721 155023 294749 155051
rect 294783 155023 294811 155051
rect 294597 154961 294625 154989
rect 294659 154961 294687 154989
rect 294721 154961 294749 154989
rect 294783 154961 294811 154989
rect 296457 239147 296485 239175
rect 296519 239147 296547 239175
rect 296581 239147 296609 239175
rect 296643 239147 296671 239175
rect 296457 239085 296485 239113
rect 296519 239085 296547 239113
rect 296581 239085 296609 239113
rect 296643 239085 296671 239113
rect 296457 239023 296485 239051
rect 296519 239023 296547 239051
rect 296581 239023 296609 239051
rect 296643 239023 296671 239051
rect 296457 238961 296485 238989
rect 296519 238961 296547 238989
rect 296581 238961 296609 238989
rect 296643 238961 296671 238989
rect 296457 230147 296485 230175
rect 296519 230147 296547 230175
rect 296581 230147 296609 230175
rect 296643 230147 296671 230175
rect 296457 230085 296485 230113
rect 296519 230085 296547 230113
rect 296581 230085 296609 230113
rect 296643 230085 296671 230113
rect 296457 230023 296485 230051
rect 296519 230023 296547 230051
rect 296581 230023 296609 230051
rect 296643 230023 296671 230051
rect 296457 229961 296485 229989
rect 296519 229961 296547 229989
rect 296581 229961 296609 229989
rect 296643 229961 296671 229989
rect 296457 221147 296485 221175
rect 296519 221147 296547 221175
rect 296581 221147 296609 221175
rect 296643 221147 296671 221175
rect 296457 221085 296485 221113
rect 296519 221085 296547 221113
rect 296581 221085 296609 221113
rect 296643 221085 296671 221113
rect 296457 221023 296485 221051
rect 296519 221023 296547 221051
rect 296581 221023 296609 221051
rect 296643 221023 296671 221051
rect 296457 220961 296485 220989
rect 296519 220961 296547 220989
rect 296581 220961 296609 220989
rect 296643 220961 296671 220989
rect 296457 212147 296485 212175
rect 296519 212147 296547 212175
rect 296581 212147 296609 212175
rect 296643 212147 296671 212175
rect 296457 212085 296485 212113
rect 296519 212085 296547 212113
rect 296581 212085 296609 212113
rect 296643 212085 296671 212113
rect 296457 212023 296485 212051
rect 296519 212023 296547 212051
rect 296581 212023 296609 212051
rect 296643 212023 296671 212051
rect 296457 211961 296485 211989
rect 296519 211961 296547 211989
rect 296581 211961 296609 211989
rect 296643 211961 296671 211989
rect 296457 203147 296485 203175
rect 296519 203147 296547 203175
rect 296581 203147 296609 203175
rect 296643 203147 296671 203175
rect 296457 203085 296485 203113
rect 296519 203085 296547 203113
rect 296581 203085 296609 203113
rect 296643 203085 296671 203113
rect 296457 203023 296485 203051
rect 296519 203023 296547 203051
rect 296581 203023 296609 203051
rect 296643 203023 296671 203051
rect 296457 202961 296485 202989
rect 296519 202961 296547 202989
rect 296581 202961 296609 202989
rect 296643 202961 296671 202989
rect 296457 194147 296485 194175
rect 296519 194147 296547 194175
rect 296581 194147 296609 194175
rect 296643 194147 296671 194175
rect 296457 194085 296485 194113
rect 296519 194085 296547 194113
rect 296581 194085 296609 194113
rect 296643 194085 296671 194113
rect 296457 194023 296485 194051
rect 296519 194023 296547 194051
rect 296581 194023 296609 194051
rect 296643 194023 296671 194051
rect 296457 193961 296485 193989
rect 296519 193961 296547 193989
rect 296581 193961 296609 193989
rect 296643 193961 296671 193989
rect 296457 185147 296485 185175
rect 296519 185147 296547 185175
rect 296581 185147 296609 185175
rect 296643 185147 296671 185175
rect 296457 185085 296485 185113
rect 296519 185085 296547 185113
rect 296581 185085 296609 185113
rect 296643 185085 296671 185113
rect 296457 185023 296485 185051
rect 296519 185023 296547 185051
rect 296581 185023 296609 185051
rect 296643 185023 296671 185051
rect 296457 184961 296485 184989
rect 296519 184961 296547 184989
rect 296581 184961 296609 184989
rect 296643 184961 296671 184989
rect 296457 176147 296485 176175
rect 296519 176147 296547 176175
rect 296581 176147 296609 176175
rect 296643 176147 296671 176175
rect 296457 176085 296485 176113
rect 296519 176085 296547 176113
rect 296581 176085 296609 176113
rect 296643 176085 296671 176113
rect 296457 176023 296485 176051
rect 296519 176023 296547 176051
rect 296581 176023 296609 176051
rect 296643 176023 296671 176051
rect 296457 175961 296485 175989
rect 296519 175961 296547 175989
rect 296581 175961 296609 175989
rect 296643 175961 296671 175989
rect 296457 167147 296485 167175
rect 296519 167147 296547 167175
rect 296581 167147 296609 167175
rect 296643 167147 296671 167175
rect 296457 167085 296485 167113
rect 296519 167085 296547 167113
rect 296581 167085 296609 167113
rect 296643 167085 296671 167113
rect 296457 167023 296485 167051
rect 296519 167023 296547 167051
rect 296581 167023 296609 167051
rect 296643 167023 296671 167051
rect 296457 166961 296485 166989
rect 296519 166961 296547 166989
rect 296581 166961 296609 166989
rect 296643 166961 296671 166989
rect 296457 158147 296485 158175
rect 296519 158147 296547 158175
rect 296581 158147 296609 158175
rect 296643 158147 296671 158175
rect 296457 158085 296485 158113
rect 296519 158085 296547 158113
rect 296581 158085 296609 158113
rect 296643 158085 296671 158113
rect 296457 158023 296485 158051
rect 296519 158023 296547 158051
rect 296581 158023 296609 158051
rect 296643 158023 296671 158051
rect 296457 157961 296485 157989
rect 296519 157961 296547 157989
rect 296581 157961 296609 157989
rect 296643 157961 296671 157989
rect 294597 146147 294625 146175
rect 294659 146147 294687 146175
rect 294721 146147 294749 146175
rect 294783 146147 294811 146175
rect 294597 146085 294625 146113
rect 294659 146085 294687 146113
rect 294721 146085 294749 146113
rect 294783 146085 294811 146113
rect 294597 146023 294625 146051
rect 294659 146023 294687 146051
rect 294721 146023 294749 146051
rect 294783 146023 294811 146051
rect 294597 145961 294625 145989
rect 294659 145961 294687 145989
rect 294721 145961 294749 145989
rect 294783 145961 294811 145989
rect 294597 137147 294625 137175
rect 294659 137147 294687 137175
rect 294721 137147 294749 137175
rect 294783 137147 294811 137175
rect 294597 137085 294625 137113
rect 294659 137085 294687 137113
rect 294721 137085 294749 137113
rect 294783 137085 294811 137113
rect 294597 137023 294625 137051
rect 294659 137023 294687 137051
rect 294721 137023 294749 137051
rect 294783 137023 294811 137051
rect 294597 136961 294625 136989
rect 294659 136961 294687 136989
rect 294721 136961 294749 136989
rect 294783 136961 294811 136989
rect 294597 128147 294625 128175
rect 294659 128147 294687 128175
rect 294721 128147 294749 128175
rect 294783 128147 294811 128175
rect 294597 128085 294625 128113
rect 294659 128085 294687 128113
rect 294721 128085 294749 128113
rect 294783 128085 294811 128113
rect 294597 128023 294625 128051
rect 294659 128023 294687 128051
rect 294721 128023 294749 128051
rect 294783 128023 294811 128051
rect 294597 127961 294625 127989
rect 294659 127961 294687 127989
rect 294721 127961 294749 127989
rect 294783 127961 294811 127989
rect 296457 149147 296485 149175
rect 296519 149147 296547 149175
rect 296581 149147 296609 149175
rect 296643 149147 296671 149175
rect 296457 149085 296485 149113
rect 296519 149085 296547 149113
rect 296581 149085 296609 149113
rect 296643 149085 296671 149113
rect 296457 149023 296485 149051
rect 296519 149023 296547 149051
rect 296581 149023 296609 149051
rect 296643 149023 296671 149051
rect 296457 148961 296485 148989
rect 296519 148961 296547 148989
rect 296581 148961 296609 148989
rect 296643 148961 296671 148989
rect 296457 140147 296485 140175
rect 296519 140147 296547 140175
rect 296581 140147 296609 140175
rect 296643 140147 296671 140175
rect 296457 140085 296485 140113
rect 296519 140085 296547 140113
rect 296581 140085 296609 140113
rect 296643 140085 296671 140113
rect 296457 140023 296485 140051
rect 296519 140023 296547 140051
rect 296581 140023 296609 140051
rect 296643 140023 296671 140051
rect 296457 139961 296485 139989
rect 296519 139961 296547 139989
rect 296581 139961 296609 139989
rect 296643 139961 296671 139989
rect 296457 131147 296485 131175
rect 296519 131147 296547 131175
rect 296581 131147 296609 131175
rect 296643 131147 296671 131175
rect 296457 131085 296485 131113
rect 296519 131085 296547 131113
rect 296581 131085 296609 131113
rect 296643 131085 296671 131113
rect 296457 131023 296485 131051
rect 296519 131023 296547 131051
rect 296581 131023 296609 131051
rect 296643 131023 296671 131051
rect 296457 130961 296485 130989
rect 296519 130961 296547 130989
rect 296581 130961 296609 130989
rect 296643 130961 296671 130989
rect 294597 119147 294625 119175
rect 294659 119147 294687 119175
rect 294721 119147 294749 119175
rect 294783 119147 294811 119175
rect 294597 119085 294625 119113
rect 294659 119085 294687 119113
rect 294721 119085 294749 119113
rect 294783 119085 294811 119113
rect 294597 119023 294625 119051
rect 294659 119023 294687 119051
rect 294721 119023 294749 119051
rect 294783 119023 294811 119051
rect 294597 118961 294625 118989
rect 294659 118961 294687 118989
rect 294721 118961 294749 118989
rect 294783 118961 294811 118989
rect 294597 110147 294625 110175
rect 294659 110147 294687 110175
rect 294721 110147 294749 110175
rect 294783 110147 294811 110175
rect 294597 110085 294625 110113
rect 294659 110085 294687 110113
rect 294721 110085 294749 110113
rect 294783 110085 294811 110113
rect 294597 110023 294625 110051
rect 294659 110023 294687 110051
rect 294721 110023 294749 110051
rect 294783 110023 294811 110051
rect 294597 109961 294625 109989
rect 294659 109961 294687 109989
rect 294721 109961 294749 109989
rect 294783 109961 294811 109989
rect 294597 101147 294625 101175
rect 294659 101147 294687 101175
rect 294721 101147 294749 101175
rect 294783 101147 294811 101175
rect 294597 101085 294625 101113
rect 294659 101085 294687 101113
rect 294721 101085 294749 101113
rect 294783 101085 294811 101113
rect 294597 101023 294625 101051
rect 294659 101023 294687 101051
rect 294721 101023 294749 101051
rect 294783 101023 294811 101051
rect 294597 100961 294625 100989
rect 294659 100961 294687 100989
rect 294721 100961 294749 100989
rect 294783 100961 294811 100989
rect 294597 92147 294625 92175
rect 294659 92147 294687 92175
rect 294721 92147 294749 92175
rect 294783 92147 294811 92175
rect 294597 92085 294625 92113
rect 294659 92085 294687 92113
rect 294721 92085 294749 92113
rect 294783 92085 294811 92113
rect 294597 92023 294625 92051
rect 294659 92023 294687 92051
rect 294721 92023 294749 92051
rect 294783 92023 294811 92051
rect 294597 91961 294625 91989
rect 294659 91961 294687 91989
rect 294721 91961 294749 91989
rect 294783 91961 294811 91989
rect 294597 83147 294625 83175
rect 294659 83147 294687 83175
rect 294721 83147 294749 83175
rect 294783 83147 294811 83175
rect 294597 83085 294625 83113
rect 294659 83085 294687 83113
rect 294721 83085 294749 83113
rect 294783 83085 294811 83113
rect 294597 83023 294625 83051
rect 294659 83023 294687 83051
rect 294721 83023 294749 83051
rect 294783 83023 294811 83051
rect 294597 82961 294625 82989
rect 294659 82961 294687 82989
rect 294721 82961 294749 82989
rect 294783 82961 294811 82989
rect 296457 122147 296485 122175
rect 296519 122147 296547 122175
rect 296581 122147 296609 122175
rect 296643 122147 296671 122175
rect 296457 122085 296485 122113
rect 296519 122085 296547 122113
rect 296581 122085 296609 122113
rect 296643 122085 296671 122113
rect 296457 122023 296485 122051
rect 296519 122023 296547 122051
rect 296581 122023 296609 122051
rect 296643 122023 296671 122051
rect 296457 121961 296485 121989
rect 296519 121961 296547 121989
rect 296581 121961 296609 121989
rect 296643 121961 296671 121989
rect 296457 113147 296485 113175
rect 296519 113147 296547 113175
rect 296581 113147 296609 113175
rect 296643 113147 296671 113175
rect 296457 113085 296485 113113
rect 296519 113085 296547 113113
rect 296581 113085 296609 113113
rect 296643 113085 296671 113113
rect 296457 113023 296485 113051
rect 296519 113023 296547 113051
rect 296581 113023 296609 113051
rect 296643 113023 296671 113051
rect 296457 112961 296485 112989
rect 296519 112961 296547 112989
rect 296581 112961 296609 112989
rect 296643 112961 296671 112989
rect 296457 104147 296485 104175
rect 296519 104147 296547 104175
rect 296581 104147 296609 104175
rect 296643 104147 296671 104175
rect 296457 104085 296485 104113
rect 296519 104085 296547 104113
rect 296581 104085 296609 104113
rect 296643 104085 296671 104113
rect 296457 104023 296485 104051
rect 296519 104023 296547 104051
rect 296581 104023 296609 104051
rect 296643 104023 296671 104051
rect 296457 103961 296485 103989
rect 296519 103961 296547 103989
rect 296581 103961 296609 103989
rect 296643 103961 296671 103989
rect 296457 95147 296485 95175
rect 296519 95147 296547 95175
rect 296581 95147 296609 95175
rect 296643 95147 296671 95175
rect 296457 95085 296485 95113
rect 296519 95085 296547 95113
rect 296581 95085 296609 95113
rect 296643 95085 296671 95113
rect 296457 95023 296485 95051
rect 296519 95023 296547 95051
rect 296581 95023 296609 95051
rect 296643 95023 296671 95051
rect 296457 94961 296485 94989
rect 296519 94961 296547 94989
rect 296581 94961 296609 94989
rect 296643 94961 296671 94989
rect 296457 86147 296485 86175
rect 296519 86147 296547 86175
rect 296581 86147 296609 86175
rect 296643 86147 296671 86175
rect 296457 86085 296485 86113
rect 296519 86085 296547 86113
rect 296581 86085 296609 86113
rect 296643 86085 296671 86113
rect 296457 86023 296485 86051
rect 296519 86023 296547 86051
rect 296581 86023 296609 86051
rect 296643 86023 296671 86051
rect 296457 85961 296485 85989
rect 296519 85961 296547 85989
rect 296581 85961 296609 85989
rect 296643 85961 296671 85989
rect 296457 77147 296485 77175
rect 296519 77147 296547 77175
rect 296581 77147 296609 77175
rect 296643 77147 296671 77175
rect 296457 77085 296485 77113
rect 296519 77085 296547 77113
rect 296581 77085 296609 77113
rect 296643 77085 296671 77113
rect 296457 77023 296485 77051
rect 296519 77023 296547 77051
rect 296581 77023 296609 77051
rect 296643 77023 296671 77051
rect 296457 76961 296485 76989
rect 296519 76961 296547 76989
rect 296581 76961 296609 76989
rect 296643 76961 296671 76989
rect 294597 74147 294625 74175
rect 294659 74147 294687 74175
rect 294721 74147 294749 74175
rect 294783 74147 294811 74175
rect 294597 74085 294625 74113
rect 294659 74085 294687 74113
rect 294721 74085 294749 74113
rect 294783 74085 294811 74113
rect 294597 74023 294625 74051
rect 294659 74023 294687 74051
rect 294721 74023 294749 74051
rect 294783 74023 294811 74051
rect 294597 73961 294625 73989
rect 294659 73961 294687 73989
rect 294721 73961 294749 73989
rect 294783 73961 294811 73989
rect 294597 65147 294625 65175
rect 294659 65147 294687 65175
rect 294721 65147 294749 65175
rect 294783 65147 294811 65175
rect 294597 65085 294625 65113
rect 294659 65085 294687 65113
rect 294721 65085 294749 65113
rect 294783 65085 294811 65113
rect 294597 65023 294625 65051
rect 294659 65023 294687 65051
rect 294721 65023 294749 65051
rect 294783 65023 294811 65051
rect 294597 64961 294625 64989
rect 294659 64961 294687 64989
rect 294721 64961 294749 64989
rect 294783 64961 294811 64989
rect 294597 56147 294625 56175
rect 294659 56147 294687 56175
rect 294721 56147 294749 56175
rect 294783 56147 294811 56175
rect 294597 56085 294625 56113
rect 294659 56085 294687 56113
rect 294721 56085 294749 56113
rect 294783 56085 294811 56113
rect 294597 56023 294625 56051
rect 294659 56023 294687 56051
rect 294721 56023 294749 56051
rect 294783 56023 294811 56051
rect 294597 55961 294625 55989
rect 294659 55961 294687 55989
rect 294721 55961 294749 55989
rect 294783 55961 294811 55989
rect 294597 47147 294625 47175
rect 294659 47147 294687 47175
rect 294721 47147 294749 47175
rect 294783 47147 294811 47175
rect 294597 47085 294625 47113
rect 294659 47085 294687 47113
rect 294721 47085 294749 47113
rect 294783 47085 294811 47113
rect 294597 47023 294625 47051
rect 294659 47023 294687 47051
rect 294721 47023 294749 47051
rect 294783 47023 294811 47051
rect 294597 46961 294625 46989
rect 294659 46961 294687 46989
rect 294721 46961 294749 46989
rect 294783 46961 294811 46989
rect 294597 38147 294625 38175
rect 294659 38147 294687 38175
rect 294721 38147 294749 38175
rect 294783 38147 294811 38175
rect 294597 38085 294625 38113
rect 294659 38085 294687 38113
rect 294721 38085 294749 38113
rect 294783 38085 294811 38113
rect 294597 38023 294625 38051
rect 294659 38023 294687 38051
rect 294721 38023 294749 38051
rect 294783 38023 294811 38051
rect 294597 37961 294625 37989
rect 294659 37961 294687 37989
rect 294721 37961 294749 37989
rect 294783 37961 294811 37989
rect 294597 29147 294625 29175
rect 294659 29147 294687 29175
rect 294721 29147 294749 29175
rect 294783 29147 294811 29175
rect 294597 29085 294625 29113
rect 294659 29085 294687 29113
rect 294721 29085 294749 29113
rect 294783 29085 294811 29113
rect 294597 29023 294625 29051
rect 294659 29023 294687 29051
rect 294721 29023 294749 29051
rect 294783 29023 294811 29051
rect 294597 28961 294625 28989
rect 294659 28961 294687 28989
rect 294721 28961 294749 28989
rect 294783 28961 294811 28989
rect 294597 20147 294625 20175
rect 294659 20147 294687 20175
rect 294721 20147 294749 20175
rect 294783 20147 294811 20175
rect 294597 20085 294625 20113
rect 294659 20085 294687 20113
rect 294721 20085 294749 20113
rect 294783 20085 294811 20113
rect 294597 20023 294625 20051
rect 294659 20023 294687 20051
rect 294721 20023 294749 20051
rect 294783 20023 294811 20051
rect 294597 19961 294625 19989
rect 294659 19961 294687 19989
rect 294721 19961 294749 19989
rect 294783 19961 294811 19989
rect 294597 11147 294625 11175
rect 294659 11147 294687 11175
rect 294721 11147 294749 11175
rect 294783 11147 294811 11175
rect 294597 11085 294625 11113
rect 294659 11085 294687 11113
rect 294721 11085 294749 11113
rect 294783 11085 294811 11113
rect 294597 11023 294625 11051
rect 294659 11023 294687 11051
rect 294721 11023 294749 11051
rect 294783 11023 294811 11051
rect 294597 10961 294625 10989
rect 294659 10961 294687 10989
rect 294721 10961 294749 10989
rect 294783 10961 294811 10989
rect 294597 2147 294625 2175
rect 294659 2147 294687 2175
rect 294721 2147 294749 2175
rect 294783 2147 294811 2175
rect 294597 2085 294625 2113
rect 294659 2085 294687 2113
rect 294721 2085 294749 2113
rect 294783 2085 294811 2113
rect 294597 2023 294625 2051
rect 294659 2023 294687 2051
rect 294721 2023 294749 2051
rect 294783 2023 294811 2051
rect 294597 1961 294625 1989
rect 294659 1961 294687 1989
rect 294721 1961 294749 1989
rect 294783 1961 294811 1989
rect 294597 -108 294625 -80
rect 294659 -108 294687 -80
rect 294721 -108 294749 -80
rect 294783 -108 294811 -80
rect 294597 -170 294625 -142
rect 294659 -170 294687 -142
rect 294721 -170 294749 -142
rect 294783 -170 294811 -142
rect 294597 -232 294625 -204
rect 294659 -232 294687 -204
rect 294721 -232 294749 -204
rect 294783 -232 294811 -204
rect 294597 -294 294625 -266
rect 294659 -294 294687 -266
rect 294721 -294 294749 -266
rect 294783 -294 294811 -266
rect 296457 68147 296485 68175
rect 296519 68147 296547 68175
rect 296581 68147 296609 68175
rect 296643 68147 296671 68175
rect 296457 68085 296485 68113
rect 296519 68085 296547 68113
rect 296581 68085 296609 68113
rect 296643 68085 296671 68113
rect 296457 68023 296485 68051
rect 296519 68023 296547 68051
rect 296581 68023 296609 68051
rect 296643 68023 296671 68051
rect 296457 67961 296485 67989
rect 296519 67961 296547 67989
rect 296581 67961 296609 67989
rect 296643 67961 296671 67989
rect 296457 59147 296485 59175
rect 296519 59147 296547 59175
rect 296581 59147 296609 59175
rect 296643 59147 296671 59175
rect 296457 59085 296485 59113
rect 296519 59085 296547 59113
rect 296581 59085 296609 59113
rect 296643 59085 296671 59113
rect 296457 59023 296485 59051
rect 296519 59023 296547 59051
rect 296581 59023 296609 59051
rect 296643 59023 296671 59051
rect 296457 58961 296485 58989
rect 296519 58961 296547 58989
rect 296581 58961 296609 58989
rect 296643 58961 296671 58989
rect 296457 50147 296485 50175
rect 296519 50147 296547 50175
rect 296581 50147 296609 50175
rect 296643 50147 296671 50175
rect 296457 50085 296485 50113
rect 296519 50085 296547 50113
rect 296581 50085 296609 50113
rect 296643 50085 296671 50113
rect 296457 50023 296485 50051
rect 296519 50023 296547 50051
rect 296581 50023 296609 50051
rect 296643 50023 296671 50051
rect 296457 49961 296485 49989
rect 296519 49961 296547 49989
rect 296581 49961 296609 49989
rect 296643 49961 296671 49989
rect 296457 41147 296485 41175
rect 296519 41147 296547 41175
rect 296581 41147 296609 41175
rect 296643 41147 296671 41175
rect 296457 41085 296485 41113
rect 296519 41085 296547 41113
rect 296581 41085 296609 41113
rect 296643 41085 296671 41113
rect 296457 41023 296485 41051
rect 296519 41023 296547 41051
rect 296581 41023 296609 41051
rect 296643 41023 296671 41051
rect 296457 40961 296485 40989
rect 296519 40961 296547 40989
rect 296581 40961 296609 40989
rect 296643 40961 296671 40989
rect 296457 32147 296485 32175
rect 296519 32147 296547 32175
rect 296581 32147 296609 32175
rect 296643 32147 296671 32175
rect 296457 32085 296485 32113
rect 296519 32085 296547 32113
rect 296581 32085 296609 32113
rect 296643 32085 296671 32113
rect 296457 32023 296485 32051
rect 296519 32023 296547 32051
rect 296581 32023 296609 32051
rect 296643 32023 296671 32051
rect 296457 31961 296485 31989
rect 296519 31961 296547 31989
rect 296581 31961 296609 31989
rect 296643 31961 296671 31989
rect 296457 23147 296485 23175
rect 296519 23147 296547 23175
rect 296581 23147 296609 23175
rect 296643 23147 296671 23175
rect 296457 23085 296485 23113
rect 296519 23085 296547 23113
rect 296581 23085 296609 23113
rect 296643 23085 296671 23113
rect 296457 23023 296485 23051
rect 296519 23023 296547 23051
rect 296581 23023 296609 23051
rect 296643 23023 296671 23051
rect 296457 22961 296485 22989
rect 296519 22961 296547 22989
rect 296581 22961 296609 22989
rect 296643 22961 296671 22989
rect 296457 14147 296485 14175
rect 296519 14147 296547 14175
rect 296581 14147 296609 14175
rect 296643 14147 296671 14175
rect 296457 14085 296485 14113
rect 296519 14085 296547 14113
rect 296581 14085 296609 14113
rect 296643 14085 296671 14113
rect 296457 14023 296485 14051
rect 296519 14023 296547 14051
rect 296581 14023 296609 14051
rect 296643 14023 296671 14051
rect 296457 13961 296485 13989
rect 296519 13961 296547 13989
rect 296581 13961 296609 13989
rect 296643 13961 296671 13989
rect 296457 5147 296485 5175
rect 296519 5147 296547 5175
rect 296581 5147 296609 5175
rect 296643 5147 296671 5175
rect 296457 5085 296485 5113
rect 296519 5085 296547 5113
rect 296581 5085 296609 5113
rect 296643 5085 296671 5113
rect 296457 5023 296485 5051
rect 296519 5023 296547 5051
rect 296581 5023 296609 5051
rect 296643 5023 296671 5051
rect 296457 4961 296485 4989
rect 296519 4961 296547 4989
rect 296581 4961 296609 4989
rect 296643 4961 296671 4989
rect 298248 298578 298276 298606
rect 298310 298578 298338 298606
rect 298372 298578 298400 298606
rect 298434 298578 298462 298606
rect 298248 298516 298276 298544
rect 298310 298516 298338 298544
rect 298372 298516 298400 298544
rect 298434 298516 298462 298544
rect 298248 298454 298276 298482
rect 298310 298454 298338 298482
rect 298372 298454 298400 298482
rect 298434 298454 298462 298482
rect 298248 298392 298276 298420
rect 298310 298392 298338 298420
rect 298372 298392 298400 298420
rect 298434 298392 298462 298420
rect 298248 290147 298276 290175
rect 298310 290147 298338 290175
rect 298372 290147 298400 290175
rect 298434 290147 298462 290175
rect 298248 290085 298276 290113
rect 298310 290085 298338 290113
rect 298372 290085 298400 290113
rect 298434 290085 298462 290113
rect 298248 290023 298276 290051
rect 298310 290023 298338 290051
rect 298372 290023 298400 290051
rect 298434 290023 298462 290051
rect 298248 289961 298276 289989
rect 298310 289961 298338 289989
rect 298372 289961 298400 289989
rect 298434 289961 298462 289989
rect 298248 281147 298276 281175
rect 298310 281147 298338 281175
rect 298372 281147 298400 281175
rect 298434 281147 298462 281175
rect 298248 281085 298276 281113
rect 298310 281085 298338 281113
rect 298372 281085 298400 281113
rect 298434 281085 298462 281113
rect 298248 281023 298276 281051
rect 298310 281023 298338 281051
rect 298372 281023 298400 281051
rect 298434 281023 298462 281051
rect 298248 280961 298276 280989
rect 298310 280961 298338 280989
rect 298372 280961 298400 280989
rect 298434 280961 298462 280989
rect 298248 272147 298276 272175
rect 298310 272147 298338 272175
rect 298372 272147 298400 272175
rect 298434 272147 298462 272175
rect 298248 272085 298276 272113
rect 298310 272085 298338 272113
rect 298372 272085 298400 272113
rect 298434 272085 298462 272113
rect 298248 272023 298276 272051
rect 298310 272023 298338 272051
rect 298372 272023 298400 272051
rect 298434 272023 298462 272051
rect 298248 271961 298276 271989
rect 298310 271961 298338 271989
rect 298372 271961 298400 271989
rect 298434 271961 298462 271989
rect 298248 263147 298276 263175
rect 298310 263147 298338 263175
rect 298372 263147 298400 263175
rect 298434 263147 298462 263175
rect 298248 263085 298276 263113
rect 298310 263085 298338 263113
rect 298372 263085 298400 263113
rect 298434 263085 298462 263113
rect 298248 263023 298276 263051
rect 298310 263023 298338 263051
rect 298372 263023 298400 263051
rect 298434 263023 298462 263051
rect 298248 262961 298276 262989
rect 298310 262961 298338 262989
rect 298372 262961 298400 262989
rect 298434 262961 298462 262989
rect 298248 254147 298276 254175
rect 298310 254147 298338 254175
rect 298372 254147 298400 254175
rect 298434 254147 298462 254175
rect 298248 254085 298276 254113
rect 298310 254085 298338 254113
rect 298372 254085 298400 254113
rect 298434 254085 298462 254113
rect 298248 254023 298276 254051
rect 298310 254023 298338 254051
rect 298372 254023 298400 254051
rect 298434 254023 298462 254051
rect 298248 253961 298276 253989
rect 298310 253961 298338 253989
rect 298372 253961 298400 253989
rect 298434 253961 298462 253989
rect 298248 245147 298276 245175
rect 298310 245147 298338 245175
rect 298372 245147 298400 245175
rect 298434 245147 298462 245175
rect 298248 245085 298276 245113
rect 298310 245085 298338 245113
rect 298372 245085 298400 245113
rect 298434 245085 298462 245113
rect 298248 245023 298276 245051
rect 298310 245023 298338 245051
rect 298372 245023 298400 245051
rect 298434 245023 298462 245051
rect 298248 244961 298276 244989
rect 298310 244961 298338 244989
rect 298372 244961 298400 244989
rect 298434 244961 298462 244989
rect 298248 236147 298276 236175
rect 298310 236147 298338 236175
rect 298372 236147 298400 236175
rect 298434 236147 298462 236175
rect 298248 236085 298276 236113
rect 298310 236085 298338 236113
rect 298372 236085 298400 236113
rect 298434 236085 298462 236113
rect 298248 236023 298276 236051
rect 298310 236023 298338 236051
rect 298372 236023 298400 236051
rect 298434 236023 298462 236051
rect 298248 235961 298276 235989
rect 298310 235961 298338 235989
rect 298372 235961 298400 235989
rect 298434 235961 298462 235989
rect 298248 227147 298276 227175
rect 298310 227147 298338 227175
rect 298372 227147 298400 227175
rect 298434 227147 298462 227175
rect 298248 227085 298276 227113
rect 298310 227085 298338 227113
rect 298372 227085 298400 227113
rect 298434 227085 298462 227113
rect 298248 227023 298276 227051
rect 298310 227023 298338 227051
rect 298372 227023 298400 227051
rect 298434 227023 298462 227051
rect 298248 226961 298276 226989
rect 298310 226961 298338 226989
rect 298372 226961 298400 226989
rect 298434 226961 298462 226989
rect 298248 218147 298276 218175
rect 298310 218147 298338 218175
rect 298372 218147 298400 218175
rect 298434 218147 298462 218175
rect 298248 218085 298276 218113
rect 298310 218085 298338 218113
rect 298372 218085 298400 218113
rect 298434 218085 298462 218113
rect 298248 218023 298276 218051
rect 298310 218023 298338 218051
rect 298372 218023 298400 218051
rect 298434 218023 298462 218051
rect 298248 217961 298276 217989
rect 298310 217961 298338 217989
rect 298372 217961 298400 217989
rect 298434 217961 298462 217989
rect 298248 209147 298276 209175
rect 298310 209147 298338 209175
rect 298372 209147 298400 209175
rect 298434 209147 298462 209175
rect 298248 209085 298276 209113
rect 298310 209085 298338 209113
rect 298372 209085 298400 209113
rect 298434 209085 298462 209113
rect 298248 209023 298276 209051
rect 298310 209023 298338 209051
rect 298372 209023 298400 209051
rect 298434 209023 298462 209051
rect 298248 208961 298276 208989
rect 298310 208961 298338 208989
rect 298372 208961 298400 208989
rect 298434 208961 298462 208989
rect 298248 200147 298276 200175
rect 298310 200147 298338 200175
rect 298372 200147 298400 200175
rect 298434 200147 298462 200175
rect 298248 200085 298276 200113
rect 298310 200085 298338 200113
rect 298372 200085 298400 200113
rect 298434 200085 298462 200113
rect 298248 200023 298276 200051
rect 298310 200023 298338 200051
rect 298372 200023 298400 200051
rect 298434 200023 298462 200051
rect 298248 199961 298276 199989
rect 298310 199961 298338 199989
rect 298372 199961 298400 199989
rect 298434 199961 298462 199989
rect 298248 191147 298276 191175
rect 298310 191147 298338 191175
rect 298372 191147 298400 191175
rect 298434 191147 298462 191175
rect 298248 191085 298276 191113
rect 298310 191085 298338 191113
rect 298372 191085 298400 191113
rect 298434 191085 298462 191113
rect 298248 191023 298276 191051
rect 298310 191023 298338 191051
rect 298372 191023 298400 191051
rect 298434 191023 298462 191051
rect 298248 190961 298276 190989
rect 298310 190961 298338 190989
rect 298372 190961 298400 190989
rect 298434 190961 298462 190989
rect 298248 182147 298276 182175
rect 298310 182147 298338 182175
rect 298372 182147 298400 182175
rect 298434 182147 298462 182175
rect 298248 182085 298276 182113
rect 298310 182085 298338 182113
rect 298372 182085 298400 182113
rect 298434 182085 298462 182113
rect 298248 182023 298276 182051
rect 298310 182023 298338 182051
rect 298372 182023 298400 182051
rect 298434 182023 298462 182051
rect 298248 181961 298276 181989
rect 298310 181961 298338 181989
rect 298372 181961 298400 181989
rect 298434 181961 298462 181989
rect 298248 173147 298276 173175
rect 298310 173147 298338 173175
rect 298372 173147 298400 173175
rect 298434 173147 298462 173175
rect 298248 173085 298276 173113
rect 298310 173085 298338 173113
rect 298372 173085 298400 173113
rect 298434 173085 298462 173113
rect 298248 173023 298276 173051
rect 298310 173023 298338 173051
rect 298372 173023 298400 173051
rect 298434 173023 298462 173051
rect 298248 172961 298276 172989
rect 298310 172961 298338 172989
rect 298372 172961 298400 172989
rect 298434 172961 298462 172989
rect 298248 164147 298276 164175
rect 298310 164147 298338 164175
rect 298372 164147 298400 164175
rect 298434 164147 298462 164175
rect 298248 164085 298276 164113
rect 298310 164085 298338 164113
rect 298372 164085 298400 164113
rect 298434 164085 298462 164113
rect 298248 164023 298276 164051
rect 298310 164023 298338 164051
rect 298372 164023 298400 164051
rect 298434 164023 298462 164051
rect 298248 163961 298276 163989
rect 298310 163961 298338 163989
rect 298372 163961 298400 163989
rect 298434 163961 298462 163989
rect 298248 155147 298276 155175
rect 298310 155147 298338 155175
rect 298372 155147 298400 155175
rect 298434 155147 298462 155175
rect 298248 155085 298276 155113
rect 298310 155085 298338 155113
rect 298372 155085 298400 155113
rect 298434 155085 298462 155113
rect 298248 155023 298276 155051
rect 298310 155023 298338 155051
rect 298372 155023 298400 155051
rect 298434 155023 298462 155051
rect 298248 154961 298276 154989
rect 298310 154961 298338 154989
rect 298372 154961 298400 154989
rect 298434 154961 298462 154989
rect 298248 146147 298276 146175
rect 298310 146147 298338 146175
rect 298372 146147 298400 146175
rect 298434 146147 298462 146175
rect 298248 146085 298276 146113
rect 298310 146085 298338 146113
rect 298372 146085 298400 146113
rect 298434 146085 298462 146113
rect 298248 146023 298276 146051
rect 298310 146023 298338 146051
rect 298372 146023 298400 146051
rect 298434 146023 298462 146051
rect 298248 145961 298276 145989
rect 298310 145961 298338 145989
rect 298372 145961 298400 145989
rect 298434 145961 298462 145989
rect 298248 137147 298276 137175
rect 298310 137147 298338 137175
rect 298372 137147 298400 137175
rect 298434 137147 298462 137175
rect 298248 137085 298276 137113
rect 298310 137085 298338 137113
rect 298372 137085 298400 137113
rect 298434 137085 298462 137113
rect 298248 137023 298276 137051
rect 298310 137023 298338 137051
rect 298372 137023 298400 137051
rect 298434 137023 298462 137051
rect 298248 136961 298276 136989
rect 298310 136961 298338 136989
rect 298372 136961 298400 136989
rect 298434 136961 298462 136989
rect 298248 128147 298276 128175
rect 298310 128147 298338 128175
rect 298372 128147 298400 128175
rect 298434 128147 298462 128175
rect 298248 128085 298276 128113
rect 298310 128085 298338 128113
rect 298372 128085 298400 128113
rect 298434 128085 298462 128113
rect 298248 128023 298276 128051
rect 298310 128023 298338 128051
rect 298372 128023 298400 128051
rect 298434 128023 298462 128051
rect 298248 127961 298276 127989
rect 298310 127961 298338 127989
rect 298372 127961 298400 127989
rect 298434 127961 298462 127989
rect 298248 119147 298276 119175
rect 298310 119147 298338 119175
rect 298372 119147 298400 119175
rect 298434 119147 298462 119175
rect 298248 119085 298276 119113
rect 298310 119085 298338 119113
rect 298372 119085 298400 119113
rect 298434 119085 298462 119113
rect 298248 119023 298276 119051
rect 298310 119023 298338 119051
rect 298372 119023 298400 119051
rect 298434 119023 298462 119051
rect 298248 118961 298276 118989
rect 298310 118961 298338 118989
rect 298372 118961 298400 118989
rect 298434 118961 298462 118989
rect 298248 110147 298276 110175
rect 298310 110147 298338 110175
rect 298372 110147 298400 110175
rect 298434 110147 298462 110175
rect 298248 110085 298276 110113
rect 298310 110085 298338 110113
rect 298372 110085 298400 110113
rect 298434 110085 298462 110113
rect 298248 110023 298276 110051
rect 298310 110023 298338 110051
rect 298372 110023 298400 110051
rect 298434 110023 298462 110051
rect 298248 109961 298276 109989
rect 298310 109961 298338 109989
rect 298372 109961 298400 109989
rect 298434 109961 298462 109989
rect 298248 101147 298276 101175
rect 298310 101147 298338 101175
rect 298372 101147 298400 101175
rect 298434 101147 298462 101175
rect 298248 101085 298276 101113
rect 298310 101085 298338 101113
rect 298372 101085 298400 101113
rect 298434 101085 298462 101113
rect 298248 101023 298276 101051
rect 298310 101023 298338 101051
rect 298372 101023 298400 101051
rect 298434 101023 298462 101051
rect 298248 100961 298276 100989
rect 298310 100961 298338 100989
rect 298372 100961 298400 100989
rect 298434 100961 298462 100989
rect 298248 92147 298276 92175
rect 298310 92147 298338 92175
rect 298372 92147 298400 92175
rect 298434 92147 298462 92175
rect 298248 92085 298276 92113
rect 298310 92085 298338 92113
rect 298372 92085 298400 92113
rect 298434 92085 298462 92113
rect 298248 92023 298276 92051
rect 298310 92023 298338 92051
rect 298372 92023 298400 92051
rect 298434 92023 298462 92051
rect 298248 91961 298276 91989
rect 298310 91961 298338 91989
rect 298372 91961 298400 91989
rect 298434 91961 298462 91989
rect 298248 83147 298276 83175
rect 298310 83147 298338 83175
rect 298372 83147 298400 83175
rect 298434 83147 298462 83175
rect 298248 83085 298276 83113
rect 298310 83085 298338 83113
rect 298372 83085 298400 83113
rect 298434 83085 298462 83113
rect 298248 83023 298276 83051
rect 298310 83023 298338 83051
rect 298372 83023 298400 83051
rect 298434 83023 298462 83051
rect 298248 82961 298276 82989
rect 298310 82961 298338 82989
rect 298372 82961 298400 82989
rect 298434 82961 298462 82989
rect 298248 74147 298276 74175
rect 298310 74147 298338 74175
rect 298372 74147 298400 74175
rect 298434 74147 298462 74175
rect 298248 74085 298276 74113
rect 298310 74085 298338 74113
rect 298372 74085 298400 74113
rect 298434 74085 298462 74113
rect 298248 74023 298276 74051
rect 298310 74023 298338 74051
rect 298372 74023 298400 74051
rect 298434 74023 298462 74051
rect 298248 73961 298276 73989
rect 298310 73961 298338 73989
rect 298372 73961 298400 73989
rect 298434 73961 298462 73989
rect 298248 65147 298276 65175
rect 298310 65147 298338 65175
rect 298372 65147 298400 65175
rect 298434 65147 298462 65175
rect 298248 65085 298276 65113
rect 298310 65085 298338 65113
rect 298372 65085 298400 65113
rect 298434 65085 298462 65113
rect 298248 65023 298276 65051
rect 298310 65023 298338 65051
rect 298372 65023 298400 65051
rect 298434 65023 298462 65051
rect 298248 64961 298276 64989
rect 298310 64961 298338 64989
rect 298372 64961 298400 64989
rect 298434 64961 298462 64989
rect 298248 56147 298276 56175
rect 298310 56147 298338 56175
rect 298372 56147 298400 56175
rect 298434 56147 298462 56175
rect 298248 56085 298276 56113
rect 298310 56085 298338 56113
rect 298372 56085 298400 56113
rect 298434 56085 298462 56113
rect 298248 56023 298276 56051
rect 298310 56023 298338 56051
rect 298372 56023 298400 56051
rect 298434 56023 298462 56051
rect 298248 55961 298276 55989
rect 298310 55961 298338 55989
rect 298372 55961 298400 55989
rect 298434 55961 298462 55989
rect 298248 47147 298276 47175
rect 298310 47147 298338 47175
rect 298372 47147 298400 47175
rect 298434 47147 298462 47175
rect 298248 47085 298276 47113
rect 298310 47085 298338 47113
rect 298372 47085 298400 47113
rect 298434 47085 298462 47113
rect 298248 47023 298276 47051
rect 298310 47023 298338 47051
rect 298372 47023 298400 47051
rect 298434 47023 298462 47051
rect 298248 46961 298276 46989
rect 298310 46961 298338 46989
rect 298372 46961 298400 46989
rect 298434 46961 298462 46989
rect 298248 38147 298276 38175
rect 298310 38147 298338 38175
rect 298372 38147 298400 38175
rect 298434 38147 298462 38175
rect 298248 38085 298276 38113
rect 298310 38085 298338 38113
rect 298372 38085 298400 38113
rect 298434 38085 298462 38113
rect 298248 38023 298276 38051
rect 298310 38023 298338 38051
rect 298372 38023 298400 38051
rect 298434 38023 298462 38051
rect 298248 37961 298276 37989
rect 298310 37961 298338 37989
rect 298372 37961 298400 37989
rect 298434 37961 298462 37989
rect 298248 29147 298276 29175
rect 298310 29147 298338 29175
rect 298372 29147 298400 29175
rect 298434 29147 298462 29175
rect 298248 29085 298276 29113
rect 298310 29085 298338 29113
rect 298372 29085 298400 29113
rect 298434 29085 298462 29113
rect 298248 29023 298276 29051
rect 298310 29023 298338 29051
rect 298372 29023 298400 29051
rect 298434 29023 298462 29051
rect 298248 28961 298276 28989
rect 298310 28961 298338 28989
rect 298372 28961 298400 28989
rect 298434 28961 298462 28989
rect 298248 20147 298276 20175
rect 298310 20147 298338 20175
rect 298372 20147 298400 20175
rect 298434 20147 298462 20175
rect 298248 20085 298276 20113
rect 298310 20085 298338 20113
rect 298372 20085 298400 20113
rect 298434 20085 298462 20113
rect 298248 20023 298276 20051
rect 298310 20023 298338 20051
rect 298372 20023 298400 20051
rect 298434 20023 298462 20051
rect 298248 19961 298276 19989
rect 298310 19961 298338 19989
rect 298372 19961 298400 19989
rect 298434 19961 298462 19989
rect 298248 11147 298276 11175
rect 298310 11147 298338 11175
rect 298372 11147 298400 11175
rect 298434 11147 298462 11175
rect 298248 11085 298276 11113
rect 298310 11085 298338 11113
rect 298372 11085 298400 11113
rect 298434 11085 298462 11113
rect 298248 11023 298276 11051
rect 298310 11023 298338 11051
rect 298372 11023 298400 11051
rect 298434 11023 298462 11051
rect 298248 10961 298276 10989
rect 298310 10961 298338 10989
rect 298372 10961 298400 10989
rect 298434 10961 298462 10989
rect 298248 2147 298276 2175
rect 298310 2147 298338 2175
rect 298372 2147 298400 2175
rect 298434 2147 298462 2175
rect 298248 2085 298276 2113
rect 298310 2085 298338 2113
rect 298372 2085 298400 2113
rect 298434 2085 298462 2113
rect 298248 2023 298276 2051
rect 298310 2023 298338 2051
rect 298372 2023 298400 2051
rect 298434 2023 298462 2051
rect 298248 1961 298276 1989
rect 298310 1961 298338 1989
rect 298372 1961 298400 1989
rect 298434 1961 298462 1989
rect 298248 -108 298276 -80
rect 298310 -108 298338 -80
rect 298372 -108 298400 -80
rect 298434 -108 298462 -80
rect 298248 -170 298276 -142
rect 298310 -170 298338 -142
rect 298372 -170 298400 -142
rect 298434 -170 298462 -142
rect 298248 -232 298276 -204
rect 298310 -232 298338 -204
rect 298372 -232 298400 -204
rect 298434 -232 298462 -204
rect 298248 -294 298276 -266
rect 298310 -294 298338 -266
rect 298372 -294 298400 -266
rect 298434 -294 298462 -266
rect 298728 293147 298756 293175
rect 298790 293147 298818 293175
rect 298852 293147 298880 293175
rect 298914 293147 298942 293175
rect 298728 293085 298756 293113
rect 298790 293085 298818 293113
rect 298852 293085 298880 293113
rect 298914 293085 298942 293113
rect 298728 293023 298756 293051
rect 298790 293023 298818 293051
rect 298852 293023 298880 293051
rect 298914 293023 298942 293051
rect 298728 292961 298756 292989
rect 298790 292961 298818 292989
rect 298852 292961 298880 292989
rect 298914 292961 298942 292989
rect 298728 284147 298756 284175
rect 298790 284147 298818 284175
rect 298852 284147 298880 284175
rect 298914 284147 298942 284175
rect 298728 284085 298756 284113
rect 298790 284085 298818 284113
rect 298852 284085 298880 284113
rect 298914 284085 298942 284113
rect 298728 284023 298756 284051
rect 298790 284023 298818 284051
rect 298852 284023 298880 284051
rect 298914 284023 298942 284051
rect 298728 283961 298756 283989
rect 298790 283961 298818 283989
rect 298852 283961 298880 283989
rect 298914 283961 298942 283989
rect 298728 275147 298756 275175
rect 298790 275147 298818 275175
rect 298852 275147 298880 275175
rect 298914 275147 298942 275175
rect 298728 275085 298756 275113
rect 298790 275085 298818 275113
rect 298852 275085 298880 275113
rect 298914 275085 298942 275113
rect 298728 275023 298756 275051
rect 298790 275023 298818 275051
rect 298852 275023 298880 275051
rect 298914 275023 298942 275051
rect 298728 274961 298756 274989
rect 298790 274961 298818 274989
rect 298852 274961 298880 274989
rect 298914 274961 298942 274989
rect 298728 266147 298756 266175
rect 298790 266147 298818 266175
rect 298852 266147 298880 266175
rect 298914 266147 298942 266175
rect 298728 266085 298756 266113
rect 298790 266085 298818 266113
rect 298852 266085 298880 266113
rect 298914 266085 298942 266113
rect 298728 266023 298756 266051
rect 298790 266023 298818 266051
rect 298852 266023 298880 266051
rect 298914 266023 298942 266051
rect 298728 265961 298756 265989
rect 298790 265961 298818 265989
rect 298852 265961 298880 265989
rect 298914 265961 298942 265989
rect 298728 257147 298756 257175
rect 298790 257147 298818 257175
rect 298852 257147 298880 257175
rect 298914 257147 298942 257175
rect 298728 257085 298756 257113
rect 298790 257085 298818 257113
rect 298852 257085 298880 257113
rect 298914 257085 298942 257113
rect 298728 257023 298756 257051
rect 298790 257023 298818 257051
rect 298852 257023 298880 257051
rect 298914 257023 298942 257051
rect 298728 256961 298756 256989
rect 298790 256961 298818 256989
rect 298852 256961 298880 256989
rect 298914 256961 298942 256989
rect 298728 248147 298756 248175
rect 298790 248147 298818 248175
rect 298852 248147 298880 248175
rect 298914 248147 298942 248175
rect 298728 248085 298756 248113
rect 298790 248085 298818 248113
rect 298852 248085 298880 248113
rect 298914 248085 298942 248113
rect 298728 248023 298756 248051
rect 298790 248023 298818 248051
rect 298852 248023 298880 248051
rect 298914 248023 298942 248051
rect 298728 247961 298756 247989
rect 298790 247961 298818 247989
rect 298852 247961 298880 247989
rect 298914 247961 298942 247989
rect 298728 239147 298756 239175
rect 298790 239147 298818 239175
rect 298852 239147 298880 239175
rect 298914 239147 298942 239175
rect 298728 239085 298756 239113
rect 298790 239085 298818 239113
rect 298852 239085 298880 239113
rect 298914 239085 298942 239113
rect 298728 239023 298756 239051
rect 298790 239023 298818 239051
rect 298852 239023 298880 239051
rect 298914 239023 298942 239051
rect 298728 238961 298756 238989
rect 298790 238961 298818 238989
rect 298852 238961 298880 238989
rect 298914 238961 298942 238989
rect 298728 230147 298756 230175
rect 298790 230147 298818 230175
rect 298852 230147 298880 230175
rect 298914 230147 298942 230175
rect 298728 230085 298756 230113
rect 298790 230085 298818 230113
rect 298852 230085 298880 230113
rect 298914 230085 298942 230113
rect 298728 230023 298756 230051
rect 298790 230023 298818 230051
rect 298852 230023 298880 230051
rect 298914 230023 298942 230051
rect 298728 229961 298756 229989
rect 298790 229961 298818 229989
rect 298852 229961 298880 229989
rect 298914 229961 298942 229989
rect 298728 221147 298756 221175
rect 298790 221147 298818 221175
rect 298852 221147 298880 221175
rect 298914 221147 298942 221175
rect 298728 221085 298756 221113
rect 298790 221085 298818 221113
rect 298852 221085 298880 221113
rect 298914 221085 298942 221113
rect 298728 221023 298756 221051
rect 298790 221023 298818 221051
rect 298852 221023 298880 221051
rect 298914 221023 298942 221051
rect 298728 220961 298756 220989
rect 298790 220961 298818 220989
rect 298852 220961 298880 220989
rect 298914 220961 298942 220989
rect 298728 212147 298756 212175
rect 298790 212147 298818 212175
rect 298852 212147 298880 212175
rect 298914 212147 298942 212175
rect 298728 212085 298756 212113
rect 298790 212085 298818 212113
rect 298852 212085 298880 212113
rect 298914 212085 298942 212113
rect 298728 212023 298756 212051
rect 298790 212023 298818 212051
rect 298852 212023 298880 212051
rect 298914 212023 298942 212051
rect 298728 211961 298756 211989
rect 298790 211961 298818 211989
rect 298852 211961 298880 211989
rect 298914 211961 298942 211989
rect 298728 203147 298756 203175
rect 298790 203147 298818 203175
rect 298852 203147 298880 203175
rect 298914 203147 298942 203175
rect 298728 203085 298756 203113
rect 298790 203085 298818 203113
rect 298852 203085 298880 203113
rect 298914 203085 298942 203113
rect 298728 203023 298756 203051
rect 298790 203023 298818 203051
rect 298852 203023 298880 203051
rect 298914 203023 298942 203051
rect 298728 202961 298756 202989
rect 298790 202961 298818 202989
rect 298852 202961 298880 202989
rect 298914 202961 298942 202989
rect 298728 194147 298756 194175
rect 298790 194147 298818 194175
rect 298852 194147 298880 194175
rect 298914 194147 298942 194175
rect 298728 194085 298756 194113
rect 298790 194085 298818 194113
rect 298852 194085 298880 194113
rect 298914 194085 298942 194113
rect 298728 194023 298756 194051
rect 298790 194023 298818 194051
rect 298852 194023 298880 194051
rect 298914 194023 298942 194051
rect 298728 193961 298756 193989
rect 298790 193961 298818 193989
rect 298852 193961 298880 193989
rect 298914 193961 298942 193989
rect 298728 185147 298756 185175
rect 298790 185147 298818 185175
rect 298852 185147 298880 185175
rect 298914 185147 298942 185175
rect 298728 185085 298756 185113
rect 298790 185085 298818 185113
rect 298852 185085 298880 185113
rect 298914 185085 298942 185113
rect 298728 185023 298756 185051
rect 298790 185023 298818 185051
rect 298852 185023 298880 185051
rect 298914 185023 298942 185051
rect 298728 184961 298756 184989
rect 298790 184961 298818 184989
rect 298852 184961 298880 184989
rect 298914 184961 298942 184989
rect 298728 176147 298756 176175
rect 298790 176147 298818 176175
rect 298852 176147 298880 176175
rect 298914 176147 298942 176175
rect 298728 176085 298756 176113
rect 298790 176085 298818 176113
rect 298852 176085 298880 176113
rect 298914 176085 298942 176113
rect 298728 176023 298756 176051
rect 298790 176023 298818 176051
rect 298852 176023 298880 176051
rect 298914 176023 298942 176051
rect 298728 175961 298756 175989
rect 298790 175961 298818 175989
rect 298852 175961 298880 175989
rect 298914 175961 298942 175989
rect 298728 167147 298756 167175
rect 298790 167147 298818 167175
rect 298852 167147 298880 167175
rect 298914 167147 298942 167175
rect 298728 167085 298756 167113
rect 298790 167085 298818 167113
rect 298852 167085 298880 167113
rect 298914 167085 298942 167113
rect 298728 167023 298756 167051
rect 298790 167023 298818 167051
rect 298852 167023 298880 167051
rect 298914 167023 298942 167051
rect 298728 166961 298756 166989
rect 298790 166961 298818 166989
rect 298852 166961 298880 166989
rect 298914 166961 298942 166989
rect 298728 158147 298756 158175
rect 298790 158147 298818 158175
rect 298852 158147 298880 158175
rect 298914 158147 298942 158175
rect 298728 158085 298756 158113
rect 298790 158085 298818 158113
rect 298852 158085 298880 158113
rect 298914 158085 298942 158113
rect 298728 158023 298756 158051
rect 298790 158023 298818 158051
rect 298852 158023 298880 158051
rect 298914 158023 298942 158051
rect 298728 157961 298756 157989
rect 298790 157961 298818 157989
rect 298852 157961 298880 157989
rect 298914 157961 298942 157989
rect 298728 149147 298756 149175
rect 298790 149147 298818 149175
rect 298852 149147 298880 149175
rect 298914 149147 298942 149175
rect 298728 149085 298756 149113
rect 298790 149085 298818 149113
rect 298852 149085 298880 149113
rect 298914 149085 298942 149113
rect 298728 149023 298756 149051
rect 298790 149023 298818 149051
rect 298852 149023 298880 149051
rect 298914 149023 298942 149051
rect 298728 148961 298756 148989
rect 298790 148961 298818 148989
rect 298852 148961 298880 148989
rect 298914 148961 298942 148989
rect 298728 140147 298756 140175
rect 298790 140147 298818 140175
rect 298852 140147 298880 140175
rect 298914 140147 298942 140175
rect 298728 140085 298756 140113
rect 298790 140085 298818 140113
rect 298852 140085 298880 140113
rect 298914 140085 298942 140113
rect 298728 140023 298756 140051
rect 298790 140023 298818 140051
rect 298852 140023 298880 140051
rect 298914 140023 298942 140051
rect 298728 139961 298756 139989
rect 298790 139961 298818 139989
rect 298852 139961 298880 139989
rect 298914 139961 298942 139989
rect 298728 131147 298756 131175
rect 298790 131147 298818 131175
rect 298852 131147 298880 131175
rect 298914 131147 298942 131175
rect 298728 131085 298756 131113
rect 298790 131085 298818 131113
rect 298852 131085 298880 131113
rect 298914 131085 298942 131113
rect 298728 131023 298756 131051
rect 298790 131023 298818 131051
rect 298852 131023 298880 131051
rect 298914 131023 298942 131051
rect 298728 130961 298756 130989
rect 298790 130961 298818 130989
rect 298852 130961 298880 130989
rect 298914 130961 298942 130989
rect 298728 122147 298756 122175
rect 298790 122147 298818 122175
rect 298852 122147 298880 122175
rect 298914 122147 298942 122175
rect 298728 122085 298756 122113
rect 298790 122085 298818 122113
rect 298852 122085 298880 122113
rect 298914 122085 298942 122113
rect 298728 122023 298756 122051
rect 298790 122023 298818 122051
rect 298852 122023 298880 122051
rect 298914 122023 298942 122051
rect 298728 121961 298756 121989
rect 298790 121961 298818 121989
rect 298852 121961 298880 121989
rect 298914 121961 298942 121989
rect 298728 113147 298756 113175
rect 298790 113147 298818 113175
rect 298852 113147 298880 113175
rect 298914 113147 298942 113175
rect 298728 113085 298756 113113
rect 298790 113085 298818 113113
rect 298852 113085 298880 113113
rect 298914 113085 298942 113113
rect 298728 113023 298756 113051
rect 298790 113023 298818 113051
rect 298852 113023 298880 113051
rect 298914 113023 298942 113051
rect 298728 112961 298756 112989
rect 298790 112961 298818 112989
rect 298852 112961 298880 112989
rect 298914 112961 298942 112989
rect 298728 104147 298756 104175
rect 298790 104147 298818 104175
rect 298852 104147 298880 104175
rect 298914 104147 298942 104175
rect 298728 104085 298756 104113
rect 298790 104085 298818 104113
rect 298852 104085 298880 104113
rect 298914 104085 298942 104113
rect 298728 104023 298756 104051
rect 298790 104023 298818 104051
rect 298852 104023 298880 104051
rect 298914 104023 298942 104051
rect 298728 103961 298756 103989
rect 298790 103961 298818 103989
rect 298852 103961 298880 103989
rect 298914 103961 298942 103989
rect 298728 95147 298756 95175
rect 298790 95147 298818 95175
rect 298852 95147 298880 95175
rect 298914 95147 298942 95175
rect 298728 95085 298756 95113
rect 298790 95085 298818 95113
rect 298852 95085 298880 95113
rect 298914 95085 298942 95113
rect 298728 95023 298756 95051
rect 298790 95023 298818 95051
rect 298852 95023 298880 95051
rect 298914 95023 298942 95051
rect 298728 94961 298756 94989
rect 298790 94961 298818 94989
rect 298852 94961 298880 94989
rect 298914 94961 298942 94989
rect 298728 86147 298756 86175
rect 298790 86147 298818 86175
rect 298852 86147 298880 86175
rect 298914 86147 298942 86175
rect 298728 86085 298756 86113
rect 298790 86085 298818 86113
rect 298852 86085 298880 86113
rect 298914 86085 298942 86113
rect 298728 86023 298756 86051
rect 298790 86023 298818 86051
rect 298852 86023 298880 86051
rect 298914 86023 298942 86051
rect 298728 85961 298756 85989
rect 298790 85961 298818 85989
rect 298852 85961 298880 85989
rect 298914 85961 298942 85989
rect 298728 77147 298756 77175
rect 298790 77147 298818 77175
rect 298852 77147 298880 77175
rect 298914 77147 298942 77175
rect 298728 77085 298756 77113
rect 298790 77085 298818 77113
rect 298852 77085 298880 77113
rect 298914 77085 298942 77113
rect 298728 77023 298756 77051
rect 298790 77023 298818 77051
rect 298852 77023 298880 77051
rect 298914 77023 298942 77051
rect 298728 76961 298756 76989
rect 298790 76961 298818 76989
rect 298852 76961 298880 76989
rect 298914 76961 298942 76989
rect 298728 68147 298756 68175
rect 298790 68147 298818 68175
rect 298852 68147 298880 68175
rect 298914 68147 298942 68175
rect 298728 68085 298756 68113
rect 298790 68085 298818 68113
rect 298852 68085 298880 68113
rect 298914 68085 298942 68113
rect 298728 68023 298756 68051
rect 298790 68023 298818 68051
rect 298852 68023 298880 68051
rect 298914 68023 298942 68051
rect 298728 67961 298756 67989
rect 298790 67961 298818 67989
rect 298852 67961 298880 67989
rect 298914 67961 298942 67989
rect 298728 59147 298756 59175
rect 298790 59147 298818 59175
rect 298852 59147 298880 59175
rect 298914 59147 298942 59175
rect 298728 59085 298756 59113
rect 298790 59085 298818 59113
rect 298852 59085 298880 59113
rect 298914 59085 298942 59113
rect 298728 59023 298756 59051
rect 298790 59023 298818 59051
rect 298852 59023 298880 59051
rect 298914 59023 298942 59051
rect 298728 58961 298756 58989
rect 298790 58961 298818 58989
rect 298852 58961 298880 58989
rect 298914 58961 298942 58989
rect 298728 50147 298756 50175
rect 298790 50147 298818 50175
rect 298852 50147 298880 50175
rect 298914 50147 298942 50175
rect 298728 50085 298756 50113
rect 298790 50085 298818 50113
rect 298852 50085 298880 50113
rect 298914 50085 298942 50113
rect 298728 50023 298756 50051
rect 298790 50023 298818 50051
rect 298852 50023 298880 50051
rect 298914 50023 298942 50051
rect 298728 49961 298756 49989
rect 298790 49961 298818 49989
rect 298852 49961 298880 49989
rect 298914 49961 298942 49989
rect 298728 41147 298756 41175
rect 298790 41147 298818 41175
rect 298852 41147 298880 41175
rect 298914 41147 298942 41175
rect 298728 41085 298756 41113
rect 298790 41085 298818 41113
rect 298852 41085 298880 41113
rect 298914 41085 298942 41113
rect 298728 41023 298756 41051
rect 298790 41023 298818 41051
rect 298852 41023 298880 41051
rect 298914 41023 298942 41051
rect 298728 40961 298756 40989
rect 298790 40961 298818 40989
rect 298852 40961 298880 40989
rect 298914 40961 298942 40989
rect 298728 32147 298756 32175
rect 298790 32147 298818 32175
rect 298852 32147 298880 32175
rect 298914 32147 298942 32175
rect 298728 32085 298756 32113
rect 298790 32085 298818 32113
rect 298852 32085 298880 32113
rect 298914 32085 298942 32113
rect 298728 32023 298756 32051
rect 298790 32023 298818 32051
rect 298852 32023 298880 32051
rect 298914 32023 298942 32051
rect 298728 31961 298756 31989
rect 298790 31961 298818 31989
rect 298852 31961 298880 31989
rect 298914 31961 298942 31989
rect 298728 23147 298756 23175
rect 298790 23147 298818 23175
rect 298852 23147 298880 23175
rect 298914 23147 298942 23175
rect 298728 23085 298756 23113
rect 298790 23085 298818 23113
rect 298852 23085 298880 23113
rect 298914 23085 298942 23113
rect 298728 23023 298756 23051
rect 298790 23023 298818 23051
rect 298852 23023 298880 23051
rect 298914 23023 298942 23051
rect 298728 22961 298756 22989
rect 298790 22961 298818 22989
rect 298852 22961 298880 22989
rect 298914 22961 298942 22989
rect 298728 14147 298756 14175
rect 298790 14147 298818 14175
rect 298852 14147 298880 14175
rect 298914 14147 298942 14175
rect 298728 14085 298756 14113
rect 298790 14085 298818 14113
rect 298852 14085 298880 14113
rect 298914 14085 298942 14113
rect 298728 14023 298756 14051
rect 298790 14023 298818 14051
rect 298852 14023 298880 14051
rect 298914 14023 298942 14051
rect 298728 13961 298756 13989
rect 298790 13961 298818 13989
rect 298852 13961 298880 13989
rect 298914 13961 298942 13989
rect 298728 5147 298756 5175
rect 298790 5147 298818 5175
rect 298852 5147 298880 5175
rect 298914 5147 298942 5175
rect 298728 5085 298756 5113
rect 298790 5085 298818 5113
rect 298852 5085 298880 5113
rect 298914 5085 298942 5113
rect 298728 5023 298756 5051
rect 298790 5023 298818 5051
rect 298852 5023 298880 5051
rect 298914 5023 298942 5051
rect 298728 4961 298756 4989
rect 298790 4961 298818 4989
rect 298852 4961 298880 4989
rect 298914 4961 298942 4989
rect 296457 -588 296485 -560
rect 296519 -588 296547 -560
rect 296581 -588 296609 -560
rect 296643 -588 296671 -560
rect 296457 -650 296485 -622
rect 296519 -650 296547 -622
rect 296581 -650 296609 -622
rect 296643 -650 296671 -622
rect 296457 -712 296485 -684
rect 296519 -712 296547 -684
rect 296581 -712 296609 -684
rect 296643 -712 296671 -684
rect 296457 -774 296485 -746
rect 296519 -774 296547 -746
rect 296581 -774 296609 -746
rect 296643 -774 296671 -746
rect 298728 -588 298756 -560
rect 298790 -588 298818 -560
rect 298852 -588 298880 -560
rect 298914 -588 298942 -560
rect 298728 -650 298756 -622
rect 298790 -650 298818 -622
rect 298852 -650 298880 -622
rect 298914 -650 298942 -622
rect 298728 -712 298756 -684
rect 298790 -712 298818 -684
rect 298852 -712 298880 -684
rect 298914 -712 298942 -684
rect 298728 -774 298756 -746
rect 298790 -774 298818 -746
rect 298852 -774 298880 -746
rect 298914 -774 298942 -746
<< metal5 >>
rect -958 299086 298990 299134
rect -958 299058 -910 299086
rect -882 299058 -848 299086
rect -820 299058 -786 299086
rect -758 299058 -724 299086
rect -696 299058 4617 299086
rect 4645 299058 4679 299086
rect 4707 299058 4741 299086
rect 4769 299058 4803 299086
rect 4831 299058 19977 299086
rect 20005 299058 20039 299086
rect 20067 299058 20101 299086
rect 20129 299058 20163 299086
rect 20191 299058 35337 299086
rect 35365 299058 35399 299086
rect 35427 299058 35461 299086
rect 35489 299058 35523 299086
rect 35551 299058 50697 299086
rect 50725 299058 50759 299086
rect 50787 299058 50821 299086
rect 50849 299058 50883 299086
rect 50911 299058 66057 299086
rect 66085 299058 66119 299086
rect 66147 299058 66181 299086
rect 66209 299058 66243 299086
rect 66271 299058 81417 299086
rect 81445 299058 81479 299086
rect 81507 299058 81541 299086
rect 81569 299058 81603 299086
rect 81631 299058 96777 299086
rect 96805 299058 96839 299086
rect 96867 299058 96901 299086
rect 96929 299058 96963 299086
rect 96991 299058 112137 299086
rect 112165 299058 112199 299086
rect 112227 299058 112261 299086
rect 112289 299058 112323 299086
rect 112351 299058 127497 299086
rect 127525 299058 127559 299086
rect 127587 299058 127621 299086
rect 127649 299058 127683 299086
rect 127711 299058 142857 299086
rect 142885 299058 142919 299086
rect 142947 299058 142981 299086
rect 143009 299058 143043 299086
rect 143071 299058 158217 299086
rect 158245 299058 158279 299086
rect 158307 299058 158341 299086
rect 158369 299058 158403 299086
rect 158431 299058 173577 299086
rect 173605 299058 173639 299086
rect 173667 299058 173701 299086
rect 173729 299058 173763 299086
rect 173791 299058 188937 299086
rect 188965 299058 188999 299086
rect 189027 299058 189061 299086
rect 189089 299058 189123 299086
rect 189151 299058 204297 299086
rect 204325 299058 204359 299086
rect 204387 299058 204421 299086
rect 204449 299058 204483 299086
rect 204511 299058 219657 299086
rect 219685 299058 219719 299086
rect 219747 299058 219781 299086
rect 219809 299058 219843 299086
rect 219871 299058 235017 299086
rect 235045 299058 235079 299086
rect 235107 299058 235141 299086
rect 235169 299058 235203 299086
rect 235231 299058 250377 299086
rect 250405 299058 250439 299086
rect 250467 299058 250501 299086
rect 250529 299058 250563 299086
rect 250591 299058 265737 299086
rect 265765 299058 265799 299086
rect 265827 299058 265861 299086
rect 265889 299058 265923 299086
rect 265951 299058 281097 299086
rect 281125 299058 281159 299086
rect 281187 299058 281221 299086
rect 281249 299058 281283 299086
rect 281311 299058 296457 299086
rect 296485 299058 296519 299086
rect 296547 299058 296581 299086
rect 296609 299058 296643 299086
rect 296671 299058 298728 299086
rect 298756 299058 298790 299086
rect 298818 299058 298852 299086
rect 298880 299058 298914 299086
rect 298942 299058 298990 299086
rect -958 299024 298990 299058
rect -958 298996 -910 299024
rect -882 298996 -848 299024
rect -820 298996 -786 299024
rect -758 298996 -724 299024
rect -696 298996 4617 299024
rect 4645 298996 4679 299024
rect 4707 298996 4741 299024
rect 4769 298996 4803 299024
rect 4831 298996 19977 299024
rect 20005 298996 20039 299024
rect 20067 298996 20101 299024
rect 20129 298996 20163 299024
rect 20191 298996 35337 299024
rect 35365 298996 35399 299024
rect 35427 298996 35461 299024
rect 35489 298996 35523 299024
rect 35551 298996 50697 299024
rect 50725 298996 50759 299024
rect 50787 298996 50821 299024
rect 50849 298996 50883 299024
rect 50911 298996 66057 299024
rect 66085 298996 66119 299024
rect 66147 298996 66181 299024
rect 66209 298996 66243 299024
rect 66271 298996 81417 299024
rect 81445 298996 81479 299024
rect 81507 298996 81541 299024
rect 81569 298996 81603 299024
rect 81631 298996 96777 299024
rect 96805 298996 96839 299024
rect 96867 298996 96901 299024
rect 96929 298996 96963 299024
rect 96991 298996 112137 299024
rect 112165 298996 112199 299024
rect 112227 298996 112261 299024
rect 112289 298996 112323 299024
rect 112351 298996 127497 299024
rect 127525 298996 127559 299024
rect 127587 298996 127621 299024
rect 127649 298996 127683 299024
rect 127711 298996 142857 299024
rect 142885 298996 142919 299024
rect 142947 298996 142981 299024
rect 143009 298996 143043 299024
rect 143071 298996 158217 299024
rect 158245 298996 158279 299024
rect 158307 298996 158341 299024
rect 158369 298996 158403 299024
rect 158431 298996 173577 299024
rect 173605 298996 173639 299024
rect 173667 298996 173701 299024
rect 173729 298996 173763 299024
rect 173791 298996 188937 299024
rect 188965 298996 188999 299024
rect 189027 298996 189061 299024
rect 189089 298996 189123 299024
rect 189151 298996 204297 299024
rect 204325 298996 204359 299024
rect 204387 298996 204421 299024
rect 204449 298996 204483 299024
rect 204511 298996 219657 299024
rect 219685 298996 219719 299024
rect 219747 298996 219781 299024
rect 219809 298996 219843 299024
rect 219871 298996 235017 299024
rect 235045 298996 235079 299024
rect 235107 298996 235141 299024
rect 235169 298996 235203 299024
rect 235231 298996 250377 299024
rect 250405 298996 250439 299024
rect 250467 298996 250501 299024
rect 250529 298996 250563 299024
rect 250591 298996 265737 299024
rect 265765 298996 265799 299024
rect 265827 298996 265861 299024
rect 265889 298996 265923 299024
rect 265951 298996 281097 299024
rect 281125 298996 281159 299024
rect 281187 298996 281221 299024
rect 281249 298996 281283 299024
rect 281311 298996 296457 299024
rect 296485 298996 296519 299024
rect 296547 298996 296581 299024
rect 296609 298996 296643 299024
rect 296671 298996 298728 299024
rect 298756 298996 298790 299024
rect 298818 298996 298852 299024
rect 298880 298996 298914 299024
rect 298942 298996 298990 299024
rect -958 298962 298990 298996
rect -958 298934 -910 298962
rect -882 298934 -848 298962
rect -820 298934 -786 298962
rect -758 298934 -724 298962
rect -696 298934 4617 298962
rect 4645 298934 4679 298962
rect 4707 298934 4741 298962
rect 4769 298934 4803 298962
rect 4831 298934 19977 298962
rect 20005 298934 20039 298962
rect 20067 298934 20101 298962
rect 20129 298934 20163 298962
rect 20191 298934 35337 298962
rect 35365 298934 35399 298962
rect 35427 298934 35461 298962
rect 35489 298934 35523 298962
rect 35551 298934 50697 298962
rect 50725 298934 50759 298962
rect 50787 298934 50821 298962
rect 50849 298934 50883 298962
rect 50911 298934 66057 298962
rect 66085 298934 66119 298962
rect 66147 298934 66181 298962
rect 66209 298934 66243 298962
rect 66271 298934 81417 298962
rect 81445 298934 81479 298962
rect 81507 298934 81541 298962
rect 81569 298934 81603 298962
rect 81631 298934 96777 298962
rect 96805 298934 96839 298962
rect 96867 298934 96901 298962
rect 96929 298934 96963 298962
rect 96991 298934 112137 298962
rect 112165 298934 112199 298962
rect 112227 298934 112261 298962
rect 112289 298934 112323 298962
rect 112351 298934 127497 298962
rect 127525 298934 127559 298962
rect 127587 298934 127621 298962
rect 127649 298934 127683 298962
rect 127711 298934 142857 298962
rect 142885 298934 142919 298962
rect 142947 298934 142981 298962
rect 143009 298934 143043 298962
rect 143071 298934 158217 298962
rect 158245 298934 158279 298962
rect 158307 298934 158341 298962
rect 158369 298934 158403 298962
rect 158431 298934 173577 298962
rect 173605 298934 173639 298962
rect 173667 298934 173701 298962
rect 173729 298934 173763 298962
rect 173791 298934 188937 298962
rect 188965 298934 188999 298962
rect 189027 298934 189061 298962
rect 189089 298934 189123 298962
rect 189151 298934 204297 298962
rect 204325 298934 204359 298962
rect 204387 298934 204421 298962
rect 204449 298934 204483 298962
rect 204511 298934 219657 298962
rect 219685 298934 219719 298962
rect 219747 298934 219781 298962
rect 219809 298934 219843 298962
rect 219871 298934 235017 298962
rect 235045 298934 235079 298962
rect 235107 298934 235141 298962
rect 235169 298934 235203 298962
rect 235231 298934 250377 298962
rect 250405 298934 250439 298962
rect 250467 298934 250501 298962
rect 250529 298934 250563 298962
rect 250591 298934 265737 298962
rect 265765 298934 265799 298962
rect 265827 298934 265861 298962
rect 265889 298934 265923 298962
rect 265951 298934 281097 298962
rect 281125 298934 281159 298962
rect 281187 298934 281221 298962
rect 281249 298934 281283 298962
rect 281311 298934 296457 298962
rect 296485 298934 296519 298962
rect 296547 298934 296581 298962
rect 296609 298934 296643 298962
rect 296671 298934 298728 298962
rect 298756 298934 298790 298962
rect 298818 298934 298852 298962
rect 298880 298934 298914 298962
rect 298942 298934 298990 298962
rect -958 298900 298990 298934
rect -958 298872 -910 298900
rect -882 298872 -848 298900
rect -820 298872 -786 298900
rect -758 298872 -724 298900
rect -696 298872 4617 298900
rect 4645 298872 4679 298900
rect 4707 298872 4741 298900
rect 4769 298872 4803 298900
rect 4831 298872 19977 298900
rect 20005 298872 20039 298900
rect 20067 298872 20101 298900
rect 20129 298872 20163 298900
rect 20191 298872 35337 298900
rect 35365 298872 35399 298900
rect 35427 298872 35461 298900
rect 35489 298872 35523 298900
rect 35551 298872 50697 298900
rect 50725 298872 50759 298900
rect 50787 298872 50821 298900
rect 50849 298872 50883 298900
rect 50911 298872 66057 298900
rect 66085 298872 66119 298900
rect 66147 298872 66181 298900
rect 66209 298872 66243 298900
rect 66271 298872 81417 298900
rect 81445 298872 81479 298900
rect 81507 298872 81541 298900
rect 81569 298872 81603 298900
rect 81631 298872 96777 298900
rect 96805 298872 96839 298900
rect 96867 298872 96901 298900
rect 96929 298872 96963 298900
rect 96991 298872 112137 298900
rect 112165 298872 112199 298900
rect 112227 298872 112261 298900
rect 112289 298872 112323 298900
rect 112351 298872 127497 298900
rect 127525 298872 127559 298900
rect 127587 298872 127621 298900
rect 127649 298872 127683 298900
rect 127711 298872 142857 298900
rect 142885 298872 142919 298900
rect 142947 298872 142981 298900
rect 143009 298872 143043 298900
rect 143071 298872 158217 298900
rect 158245 298872 158279 298900
rect 158307 298872 158341 298900
rect 158369 298872 158403 298900
rect 158431 298872 173577 298900
rect 173605 298872 173639 298900
rect 173667 298872 173701 298900
rect 173729 298872 173763 298900
rect 173791 298872 188937 298900
rect 188965 298872 188999 298900
rect 189027 298872 189061 298900
rect 189089 298872 189123 298900
rect 189151 298872 204297 298900
rect 204325 298872 204359 298900
rect 204387 298872 204421 298900
rect 204449 298872 204483 298900
rect 204511 298872 219657 298900
rect 219685 298872 219719 298900
rect 219747 298872 219781 298900
rect 219809 298872 219843 298900
rect 219871 298872 235017 298900
rect 235045 298872 235079 298900
rect 235107 298872 235141 298900
rect 235169 298872 235203 298900
rect 235231 298872 250377 298900
rect 250405 298872 250439 298900
rect 250467 298872 250501 298900
rect 250529 298872 250563 298900
rect 250591 298872 265737 298900
rect 265765 298872 265799 298900
rect 265827 298872 265861 298900
rect 265889 298872 265923 298900
rect 265951 298872 281097 298900
rect 281125 298872 281159 298900
rect 281187 298872 281221 298900
rect 281249 298872 281283 298900
rect 281311 298872 296457 298900
rect 296485 298872 296519 298900
rect 296547 298872 296581 298900
rect 296609 298872 296643 298900
rect 296671 298872 298728 298900
rect 298756 298872 298790 298900
rect 298818 298872 298852 298900
rect 298880 298872 298914 298900
rect 298942 298872 298990 298900
rect -958 298824 298990 298872
rect -478 298606 298510 298654
rect -478 298578 -430 298606
rect -402 298578 -368 298606
rect -340 298578 -306 298606
rect -278 298578 -244 298606
rect -216 298578 2757 298606
rect 2785 298578 2819 298606
rect 2847 298578 2881 298606
rect 2909 298578 2943 298606
rect 2971 298578 18117 298606
rect 18145 298578 18179 298606
rect 18207 298578 18241 298606
rect 18269 298578 18303 298606
rect 18331 298578 33477 298606
rect 33505 298578 33539 298606
rect 33567 298578 33601 298606
rect 33629 298578 33663 298606
rect 33691 298578 48837 298606
rect 48865 298578 48899 298606
rect 48927 298578 48961 298606
rect 48989 298578 49023 298606
rect 49051 298578 64197 298606
rect 64225 298578 64259 298606
rect 64287 298578 64321 298606
rect 64349 298578 64383 298606
rect 64411 298578 79557 298606
rect 79585 298578 79619 298606
rect 79647 298578 79681 298606
rect 79709 298578 79743 298606
rect 79771 298578 94917 298606
rect 94945 298578 94979 298606
rect 95007 298578 95041 298606
rect 95069 298578 95103 298606
rect 95131 298578 110277 298606
rect 110305 298578 110339 298606
rect 110367 298578 110401 298606
rect 110429 298578 110463 298606
rect 110491 298578 125637 298606
rect 125665 298578 125699 298606
rect 125727 298578 125761 298606
rect 125789 298578 125823 298606
rect 125851 298578 140997 298606
rect 141025 298578 141059 298606
rect 141087 298578 141121 298606
rect 141149 298578 141183 298606
rect 141211 298578 156357 298606
rect 156385 298578 156419 298606
rect 156447 298578 156481 298606
rect 156509 298578 156543 298606
rect 156571 298578 171717 298606
rect 171745 298578 171779 298606
rect 171807 298578 171841 298606
rect 171869 298578 171903 298606
rect 171931 298578 187077 298606
rect 187105 298578 187139 298606
rect 187167 298578 187201 298606
rect 187229 298578 187263 298606
rect 187291 298578 202437 298606
rect 202465 298578 202499 298606
rect 202527 298578 202561 298606
rect 202589 298578 202623 298606
rect 202651 298578 217797 298606
rect 217825 298578 217859 298606
rect 217887 298578 217921 298606
rect 217949 298578 217983 298606
rect 218011 298578 233157 298606
rect 233185 298578 233219 298606
rect 233247 298578 233281 298606
rect 233309 298578 233343 298606
rect 233371 298578 248517 298606
rect 248545 298578 248579 298606
rect 248607 298578 248641 298606
rect 248669 298578 248703 298606
rect 248731 298578 263877 298606
rect 263905 298578 263939 298606
rect 263967 298578 264001 298606
rect 264029 298578 264063 298606
rect 264091 298578 279237 298606
rect 279265 298578 279299 298606
rect 279327 298578 279361 298606
rect 279389 298578 279423 298606
rect 279451 298578 294597 298606
rect 294625 298578 294659 298606
rect 294687 298578 294721 298606
rect 294749 298578 294783 298606
rect 294811 298578 298248 298606
rect 298276 298578 298310 298606
rect 298338 298578 298372 298606
rect 298400 298578 298434 298606
rect 298462 298578 298510 298606
rect -478 298544 298510 298578
rect -478 298516 -430 298544
rect -402 298516 -368 298544
rect -340 298516 -306 298544
rect -278 298516 -244 298544
rect -216 298516 2757 298544
rect 2785 298516 2819 298544
rect 2847 298516 2881 298544
rect 2909 298516 2943 298544
rect 2971 298516 18117 298544
rect 18145 298516 18179 298544
rect 18207 298516 18241 298544
rect 18269 298516 18303 298544
rect 18331 298516 33477 298544
rect 33505 298516 33539 298544
rect 33567 298516 33601 298544
rect 33629 298516 33663 298544
rect 33691 298516 48837 298544
rect 48865 298516 48899 298544
rect 48927 298516 48961 298544
rect 48989 298516 49023 298544
rect 49051 298516 64197 298544
rect 64225 298516 64259 298544
rect 64287 298516 64321 298544
rect 64349 298516 64383 298544
rect 64411 298516 79557 298544
rect 79585 298516 79619 298544
rect 79647 298516 79681 298544
rect 79709 298516 79743 298544
rect 79771 298516 94917 298544
rect 94945 298516 94979 298544
rect 95007 298516 95041 298544
rect 95069 298516 95103 298544
rect 95131 298516 110277 298544
rect 110305 298516 110339 298544
rect 110367 298516 110401 298544
rect 110429 298516 110463 298544
rect 110491 298516 125637 298544
rect 125665 298516 125699 298544
rect 125727 298516 125761 298544
rect 125789 298516 125823 298544
rect 125851 298516 140997 298544
rect 141025 298516 141059 298544
rect 141087 298516 141121 298544
rect 141149 298516 141183 298544
rect 141211 298516 156357 298544
rect 156385 298516 156419 298544
rect 156447 298516 156481 298544
rect 156509 298516 156543 298544
rect 156571 298516 171717 298544
rect 171745 298516 171779 298544
rect 171807 298516 171841 298544
rect 171869 298516 171903 298544
rect 171931 298516 187077 298544
rect 187105 298516 187139 298544
rect 187167 298516 187201 298544
rect 187229 298516 187263 298544
rect 187291 298516 202437 298544
rect 202465 298516 202499 298544
rect 202527 298516 202561 298544
rect 202589 298516 202623 298544
rect 202651 298516 217797 298544
rect 217825 298516 217859 298544
rect 217887 298516 217921 298544
rect 217949 298516 217983 298544
rect 218011 298516 233157 298544
rect 233185 298516 233219 298544
rect 233247 298516 233281 298544
rect 233309 298516 233343 298544
rect 233371 298516 248517 298544
rect 248545 298516 248579 298544
rect 248607 298516 248641 298544
rect 248669 298516 248703 298544
rect 248731 298516 263877 298544
rect 263905 298516 263939 298544
rect 263967 298516 264001 298544
rect 264029 298516 264063 298544
rect 264091 298516 279237 298544
rect 279265 298516 279299 298544
rect 279327 298516 279361 298544
rect 279389 298516 279423 298544
rect 279451 298516 294597 298544
rect 294625 298516 294659 298544
rect 294687 298516 294721 298544
rect 294749 298516 294783 298544
rect 294811 298516 298248 298544
rect 298276 298516 298310 298544
rect 298338 298516 298372 298544
rect 298400 298516 298434 298544
rect 298462 298516 298510 298544
rect -478 298482 298510 298516
rect -478 298454 -430 298482
rect -402 298454 -368 298482
rect -340 298454 -306 298482
rect -278 298454 -244 298482
rect -216 298454 2757 298482
rect 2785 298454 2819 298482
rect 2847 298454 2881 298482
rect 2909 298454 2943 298482
rect 2971 298454 18117 298482
rect 18145 298454 18179 298482
rect 18207 298454 18241 298482
rect 18269 298454 18303 298482
rect 18331 298454 33477 298482
rect 33505 298454 33539 298482
rect 33567 298454 33601 298482
rect 33629 298454 33663 298482
rect 33691 298454 48837 298482
rect 48865 298454 48899 298482
rect 48927 298454 48961 298482
rect 48989 298454 49023 298482
rect 49051 298454 64197 298482
rect 64225 298454 64259 298482
rect 64287 298454 64321 298482
rect 64349 298454 64383 298482
rect 64411 298454 79557 298482
rect 79585 298454 79619 298482
rect 79647 298454 79681 298482
rect 79709 298454 79743 298482
rect 79771 298454 94917 298482
rect 94945 298454 94979 298482
rect 95007 298454 95041 298482
rect 95069 298454 95103 298482
rect 95131 298454 110277 298482
rect 110305 298454 110339 298482
rect 110367 298454 110401 298482
rect 110429 298454 110463 298482
rect 110491 298454 125637 298482
rect 125665 298454 125699 298482
rect 125727 298454 125761 298482
rect 125789 298454 125823 298482
rect 125851 298454 140997 298482
rect 141025 298454 141059 298482
rect 141087 298454 141121 298482
rect 141149 298454 141183 298482
rect 141211 298454 156357 298482
rect 156385 298454 156419 298482
rect 156447 298454 156481 298482
rect 156509 298454 156543 298482
rect 156571 298454 171717 298482
rect 171745 298454 171779 298482
rect 171807 298454 171841 298482
rect 171869 298454 171903 298482
rect 171931 298454 187077 298482
rect 187105 298454 187139 298482
rect 187167 298454 187201 298482
rect 187229 298454 187263 298482
rect 187291 298454 202437 298482
rect 202465 298454 202499 298482
rect 202527 298454 202561 298482
rect 202589 298454 202623 298482
rect 202651 298454 217797 298482
rect 217825 298454 217859 298482
rect 217887 298454 217921 298482
rect 217949 298454 217983 298482
rect 218011 298454 233157 298482
rect 233185 298454 233219 298482
rect 233247 298454 233281 298482
rect 233309 298454 233343 298482
rect 233371 298454 248517 298482
rect 248545 298454 248579 298482
rect 248607 298454 248641 298482
rect 248669 298454 248703 298482
rect 248731 298454 263877 298482
rect 263905 298454 263939 298482
rect 263967 298454 264001 298482
rect 264029 298454 264063 298482
rect 264091 298454 279237 298482
rect 279265 298454 279299 298482
rect 279327 298454 279361 298482
rect 279389 298454 279423 298482
rect 279451 298454 294597 298482
rect 294625 298454 294659 298482
rect 294687 298454 294721 298482
rect 294749 298454 294783 298482
rect 294811 298454 298248 298482
rect 298276 298454 298310 298482
rect 298338 298454 298372 298482
rect 298400 298454 298434 298482
rect 298462 298454 298510 298482
rect -478 298420 298510 298454
rect -478 298392 -430 298420
rect -402 298392 -368 298420
rect -340 298392 -306 298420
rect -278 298392 -244 298420
rect -216 298392 2757 298420
rect 2785 298392 2819 298420
rect 2847 298392 2881 298420
rect 2909 298392 2943 298420
rect 2971 298392 18117 298420
rect 18145 298392 18179 298420
rect 18207 298392 18241 298420
rect 18269 298392 18303 298420
rect 18331 298392 33477 298420
rect 33505 298392 33539 298420
rect 33567 298392 33601 298420
rect 33629 298392 33663 298420
rect 33691 298392 48837 298420
rect 48865 298392 48899 298420
rect 48927 298392 48961 298420
rect 48989 298392 49023 298420
rect 49051 298392 64197 298420
rect 64225 298392 64259 298420
rect 64287 298392 64321 298420
rect 64349 298392 64383 298420
rect 64411 298392 79557 298420
rect 79585 298392 79619 298420
rect 79647 298392 79681 298420
rect 79709 298392 79743 298420
rect 79771 298392 94917 298420
rect 94945 298392 94979 298420
rect 95007 298392 95041 298420
rect 95069 298392 95103 298420
rect 95131 298392 110277 298420
rect 110305 298392 110339 298420
rect 110367 298392 110401 298420
rect 110429 298392 110463 298420
rect 110491 298392 125637 298420
rect 125665 298392 125699 298420
rect 125727 298392 125761 298420
rect 125789 298392 125823 298420
rect 125851 298392 140997 298420
rect 141025 298392 141059 298420
rect 141087 298392 141121 298420
rect 141149 298392 141183 298420
rect 141211 298392 156357 298420
rect 156385 298392 156419 298420
rect 156447 298392 156481 298420
rect 156509 298392 156543 298420
rect 156571 298392 171717 298420
rect 171745 298392 171779 298420
rect 171807 298392 171841 298420
rect 171869 298392 171903 298420
rect 171931 298392 187077 298420
rect 187105 298392 187139 298420
rect 187167 298392 187201 298420
rect 187229 298392 187263 298420
rect 187291 298392 202437 298420
rect 202465 298392 202499 298420
rect 202527 298392 202561 298420
rect 202589 298392 202623 298420
rect 202651 298392 217797 298420
rect 217825 298392 217859 298420
rect 217887 298392 217921 298420
rect 217949 298392 217983 298420
rect 218011 298392 233157 298420
rect 233185 298392 233219 298420
rect 233247 298392 233281 298420
rect 233309 298392 233343 298420
rect 233371 298392 248517 298420
rect 248545 298392 248579 298420
rect 248607 298392 248641 298420
rect 248669 298392 248703 298420
rect 248731 298392 263877 298420
rect 263905 298392 263939 298420
rect 263967 298392 264001 298420
rect 264029 298392 264063 298420
rect 264091 298392 279237 298420
rect 279265 298392 279299 298420
rect 279327 298392 279361 298420
rect 279389 298392 279423 298420
rect 279451 298392 294597 298420
rect 294625 298392 294659 298420
rect 294687 298392 294721 298420
rect 294749 298392 294783 298420
rect 294811 298392 298248 298420
rect 298276 298392 298310 298420
rect 298338 298392 298372 298420
rect 298400 298392 298434 298420
rect 298462 298392 298510 298420
rect -478 298344 298510 298392
rect -958 293175 298990 293223
rect -958 293147 -910 293175
rect -882 293147 -848 293175
rect -820 293147 -786 293175
rect -758 293147 -724 293175
rect -696 293147 4617 293175
rect 4645 293147 4679 293175
rect 4707 293147 4741 293175
rect 4769 293147 4803 293175
rect 4831 293147 19977 293175
rect 20005 293147 20039 293175
rect 20067 293147 20101 293175
rect 20129 293147 20163 293175
rect 20191 293147 35337 293175
rect 35365 293147 35399 293175
rect 35427 293147 35461 293175
rect 35489 293147 35523 293175
rect 35551 293147 50697 293175
rect 50725 293147 50759 293175
rect 50787 293147 50821 293175
rect 50849 293147 50883 293175
rect 50911 293147 66057 293175
rect 66085 293147 66119 293175
rect 66147 293147 66181 293175
rect 66209 293147 66243 293175
rect 66271 293147 81417 293175
rect 81445 293147 81479 293175
rect 81507 293147 81541 293175
rect 81569 293147 81603 293175
rect 81631 293147 96777 293175
rect 96805 293147 96839 293175
rect 96867 293147 96901 293175
rect 96929 293147 96963 293175
rect 96991 293147 112137 293175
rect 112165 293147 112199 293175
rect 112227 293147 112261 293175
rect 112289 293147 112323 293175
rect 112351 293147 127497 293175
rect 127525 293147 127559 293175
rect 127587 293147 127621 293175
rect 127649 293147 127683 293175
rect 127711 293147 142857 293175
rect 142885 293147 142919 293175
rect 142947 293147 142981 293175
rect 143009 293147 143043 293175
rect 143071 293147 158217 293175
rect 158245 293147 158279 293175
rect 158307 293147 158341 293175
rect 158369 293147 158403 293175
rect 158431 293147 173577 293175
rect 173605 293147 173639 293175
rect 173667 293147 173701 293175
rect 173729 293147 173763 293175
rect 173791 293147 188937 293175
rect 188965 293147 188999 293175
rect 189027 293147 189061 293175
rect 189089 293147 189123 293175
rect 189151 293147 204297 293175
rect 204325 293147 204359 293175
rect 204387 293147 204421 293175
rect 204449 293147 204483 293175
rect 204511 293147 219657 293175
rect 219685 293147 219719 293175
rect 219747 293147 219781 293175
rect 219809 293147 219843 293175
rect 219871 293147 235017 293175
rect 235045 293147 235079 293175
rect 235107 293147 235141 293175
rect 235169 293147 235203 293175
rect 235231 293147 250377 293175
rect 250405 293147 250439 293175
rect 250467 293147 250501 293175
rect 250529 293147 250563 293175
rect 250591 293147 265737 293175
rect 265765 293147 265799 293175
rect 265827 293147 265861 293175
rect 265889 293147 265923 293175
rect 265951 293147 281097 293175
rect 281125 293147 281159 293175
rect 281187 293147 281221 293175
rect 281249 293147 281283 293175
rect 281311 293147 296457 293175
rect 296485 293147 296519 293175
rect 296547 293147 296581 293175
rect 296609 293147 296643 293175
rect 296671 293147 298728 293175
rect 298756 293147 298790 293175
rect 298818 293147 298852 293175
rect 298880 293147 298914 293175
rect 298942 293147 298990 293175
rect -958 293113 298990 293147
rect -958 293085 -910 293113
rect -882 293085 -848 293113
rect -820 293085 -786 293113
rect -758 293085 -724 293113
rect -696 293085 4617 293113
rect 4645 293085 4679 293113
rect 4707 293085 4741 293113
rect 4769 293085 4803 293113
rect 4831 293085 19977 293113
rect 20005 293085 20039 293113
rect 20067 293085 20101 293113
rect 20129 293085 20163 293113
rect 20191 293085 35337 293113
rect 35365 293085 35399 293113
rect 35427 293085 35461 293113
rect 35489 293085 35523 293113
rect 35551 293085 50697 293113
rect 50725 293085 50759 293113
rect 50787 293085 50821 293113
rect 50849 293085 50883 293113
rect 50911 293085 66057 293113
rect 66085 293085 66119 293113
rect 66147 293085 66181 293113
rect 66209 293085 66243 293113
rect 66271 293085 81417 293113
rect 81445 293085 81479 293113
rect 81507 293085 81541 293113
rect 81569 293085 81603 293113
rect 81631 293085 96777 293113
rect 96805 293085 96839 293113
rect 96867 293085 96901 293113
rect 96929 293085 96963 293113
rect 96991 293085 112137 293113
rect 112165 293085 112199 293113
rect 112227 293085 112261 293113
rect 112289 293085 112323 293113
rect 112351 293085 127497 293113
rect 127525 293085 127559 293113
rect 127587 293085 127621 293113
rect 127649 293085 127683 293113
rect 127711 293085 142857 293113
rect 142885 293085 142919 293113
rect 142947 293085 142981 293113
rect 143009 293085 143043 293113
rect 143071 293085 158217 293113
rect 158245 293085 158279 293113
rect 158307 293085 158341 293113
rect 158369 293085 158403 293113
rect 158431 293085 173577 293113
rect 173605 293085 173639 293113
rect 173667 293085 173701 293113
rect 173729 293085 173763 293113
rect 173791 293085 188937 293113
rect 188965 293085 188999 293113
rect 189027 293085 189061 293113
rect 189089 293085 189123 293113
rect 189151 293085 204297 293113
rect 204325 293085 204359 293113
rect 204387 293085 204421 293113
rect 204449 293085 204483 293113
rect 204511 293085 219657 293113
rect 219685 293085 219719 293113
rect 219747 293085 219781 293113
rect 219809 293085 219843 293113
rect 219871 293085 235017 293113
rect 235045 293085 235079 293113
rect 235107 293085 235141 293113
rect 235169 293085 235203 293113
rect 235231 293085 250377 293113
rect 250405 293085 250439 293113
rect 250467 293085 250501 293113
rect 250529 293085 250563 293113
rect 250591 293085 265737 293113
rect 265765 293085 265799 293113
rect 265827 293085 265861 293113
rect 265889 293085 265923 293113
rect 265951 293085 281097 293113
rect 281125 293085 281159 293113
rect 281187 293085 281221 293113
rect 281249 293085 281283 293113
rect 281311 293085 296457 293113
rect 296485 293085 296519 293113
rect 296547 293085 296581 293113
rect 296609 293085 296643 293113
rect 296671 293085 298728 293113
rect 298756 293085 298790 293113
rect 298818 293085 298852 293113
rect 298880 293085 298914 293113
rect 298942 293085 298990 293113
rect -958 293051 298990 293085
rect -958 293023 -910 293051
rect -882 293023 -848 293051
rect -820 293023 -786 293051
rect -758 293023 -724 293051
rect -696 293023 4617 293051
rect 4645 293023 4679 293051
rect 4707 293023 4741 293051
rect 4769 293023 4803 293051
rect 4831 293023 19977 293051
rect 20005 293023 20039 293051
rect 20067 293023 20101 293051
rect 20129 293023 20163 293051
rect 20191 293023 35337 293051
rect 35365 293023 35399 293051
rect 35427 293023 35461 293051
rect 35489 293023 35523 293051
rect 35551 293023 50697 293051
rect 50725 293023 50759 293051
rect 50787 293023 50821 293051
rect 50849 293023 50883 293051
rect 50911 293023 66057 293051
rect 66085 293023 66119 293051
rect 66147 293023 66181 293051
rect 66209 293023 66243 293051
rect 66271 293023 81417 293051
rect 81445 293023 81479 293051
rect 81507 293023 81541 293051
rect 81569 293023 81603 293051
rect 81631 293023 96777 293051
rect 96805 293023 96839 293051
rect 96867 293023 96901 293051
rect 96929 293023 96963 293051
rect 96991 293023 112137 293051
rect 112165 293023 112199 293051
rect 112227 293023 112261 293051
rect 112289 293023 112323 293051
rect 112351 293023 127497 293051
rect 127525 293023 127559 293051
rect 127587 293023 127621 293051
rect 127649 293023 127683 293051
rect 127711 293023 142857 293051
rect 142885 293023 142919 293051
rect 142947 293023 142981 293051
rect 143009 293023 143043 293051
rect 143071 293023 158217 293051
rect 158245 293023 158279 293051
rect 158307 293023 158341 293051
rect 158369 293023 158403 293051
rect 158431 293023 173577 293051
rect 173605 293023 173639 293051
rect 173667 293023 173701 293051
rect 173729 293023 173763 293051
rect 173791 293023 188937 293051
rect 188965 293023 188999 293051
rect 189027 293023 189061 293051
rect 189089 293023 189123 293051
rect 189151 293023 204297 293051
rect 204325 293023 204359 293051
rect 204387 293023 204421 293051
rect 204449 293023 204483 293051
rect 204511 293023 219657 293051
rect 219685 293023 219719 293051
rect 219747 293023 219781 293051
rect 219809 293023 219843 293051
rect 219871 293023 235017 293051
rect 235045 293023 235079 293051
rect 235107 293023 235141 293051
rect 235169 293023 235203 293051
rect 235231 293023 250377 293051
rect 250405 293023 250439 293051
rect 250467 293023 250501 293051
rect 250529 293023 250563 293051
rect 250591 293023 265737 293051
rect 265765 293023 265799 293051
rect 265827 293023 265861 293051
rect 265889 293023 265923 293051
rect 265951 293023 281097 293051
rect 281125 293023 281159 293051
rect 281187 293023 281221 293051
rect 281249 293023 281283 293051
rect 281311 293023 296457 293051
rect 296485 293023 296519 293051
rect 296547 293023 296581 293051
rect 296609 293023 296643 293051
rect 296671 293023 298728 293051
rect 298756 293023 298790 293051
rect 298818 293023 298852 293051
rect 298880 293023 298914 293051
rect 298942 293023 298990 293051
rect -958 292989 298990 293023
rect -958 292961 -910 292989
rect -882 292961 -848 292989
rect -820 292961 -786 292989
rect -758 292961 -724 292989
rect -696 292961 4617 292989
rect 4645 292961 4679 292989
rect 4707 292961 4741 292989
rect 4769 292961 4803 292989
rect 4831 292961 19977 292989
rect 20005 292961 20039 292989
rect 20067 292961 20101 292989
rect 20129 292961 20163 292989
rect 20191 292961 35337 292989
rect 35365 292961 35399 292989
rect 35427 292961 35461 292989
rect 35489 292961 35523 292989
rect 35551 292961 50697 292989
rect 50725 292961 50759 292989
rect 50787 292961 50821 292989
rect 50849 292961 50883 292989
rect 50911 292961 66057 292989
rect 66085 292961 66119 292989
rect 66147 292961 66181 292989
rect 66209 292961 66243 292989
rect 66271 292961 81417 292989
rect 81445 292961 81479 292989
rect 81507 292961 81541 292989
rect 81569 292961 81603 292989
rect 81631 292961 96777 292989
rect 96805 292961 96839 292989
rect 96867 292961 96901 292989
rect 96929 292961 96963 292989
rect 96991 292961 112137 292989
rect 112165 292961 112199 292989
rect 112227 292961 112261 292989
rect 112289 292961 112323 292989
rect 112351 292961 127497 292989
rect 127525 292961 127559 292989
rect 127587 292961 127621 292989
rect 127649 292961 127683 292989
rect 127711 292961 142857 292989
rect 142885 292961 142919 292989
rect 142947 292961 142981 292989
rect 143009 292961 143043 292989
rect 143071 292961 158217 292989
rect 158245 292961 158279 292989
rect 158307 292961 158341 292989
rect 158369 292961 158403 292989
rect 158431 292961 173577 292989
rect 173605 292961 173639 292989
rect 173667 292961 173701 292989
rect 173729 292961 173763 292989
rect 173791 292961 188937 292989
rect 188965 292961 188999 292989
rect 189027 292961 189061 292989
rect 189089 292961 189123 292989
rect 189151 292961 204297 292989
rect 204325 292961 204359 292989
rect 204387 292961 204421 292989
rect 204449 292961 204483 292989
rect 204511 292961 219657 292989
rect 219685 292961 219719 292989
rect 219747 292961 219781 292989
rect 219809 292961 219843 292989
rect 219871 292961 235017 292989
rect 235045 292961 235079 292989
rect 235107 292961 235141 292989
rect 235169 292961 235203 292989
rect 235231 292961 250377 292989
rect 250405 292961 250439 292989
rect 250467 292961 250501 292989
rect 250529 292961 250563 292989
rect 250591 292961 265737 292989
rect 265765 292961 265799 292989
rect 265827 292961 265861 292989
rect 265889 292961 265923 292989
rect 265951 292961 281097 292989
rect 281125 292961 281159 292989
rect 281187 292961 281221 292989
rect 281249 292961 281283 292989
rect 281311 292961 296457 292989
rect 296485 292961 296519 292989
rect 296547 292961 296581 292989
rect 296609 292961 296643 292989
rect 296671 292961 298728 292989
rect 298756 292961 298790 292989
rect 298818 292961 298852 292989
rect 298880 292961 298914 292989
rect 298942 292961 298990 292989
rect -958 292913 298990 292961
rect -958 290175 298990 290223
rect -958 290147 -430 290175
rect -402 290147 -368 290175
rect -340 290147 -306 290175
rect -278 290147 -244 290175
rect -216 290147 2757 290175
rect 2785 290147 2819 290175
rect 2847 290147 2881 290175
rect 2909 290147 2943 290175
rect 2971 290147 18117 290175
rect 18145 290147 18179 290175
rect 18207 290147 18241 290175
rect 18269 290147 18303 290175
rect 18331 290147 33477 290175
rect 33505 290147 33539 290175
rect 33567 290147 33601 290175
rect 33629 290147 33663 290175
rect 33691 290147 48837 290175
rect 48865 290147 48899 290175
rect 48927 290147 48961 290175
rect 48989 290147 49023 290175
rect 49051 290147 64197 290175
rect 64225 290147 64259 290175
rect 64287 290147 64321 290175
rect 64349 290147 64383 290175
rect 64411 290147 79557 290175
rect 79585 290147 79619 290175
rect 79647 290147 79681 290175
rect 79709 290147 79743 290175
rect 79771 290147 94917 290175
rect 94945 290147 94979 290175
rect 95007 290147 95041 290175
rect 95069 290147 95103 290175
rect 95131 290147 110277 290175
rect 110305 290147 110339 290175
rect 110367 290147 110401 290175
rect 110429 290147 110463 290175
rect 110491 290147 125637 290175
rect 125665 290147 125699 290175
rect 125727 290147 125761 290175
rect 125789 290147 125823 290175
rect 125851 290147 140997 290175
rect 141025 290147 141059 290175
rect 141087 290147 141121 290175
rect 141149 290147 141183 290175
rect 141211 290147 156357 290175
rect 156385 290147 156419 290175
rect 156447 290147 156481 290175
rect 156509 290147 156543 290175
rect 156571 290147 171717 290175
rect 171745 290147 171779 290175
rect 171807 290147 171841 290175
rect 171869 290147 171903 290175
rect 171931 290147 187077 290175
rect 187105 290147 187139 290175
rect 187167 290147 187201 290175
rect 187229 290147 187263 290175
rect 187291 290147 202437 290175
rect 202465 290147 202499 290175
rect 202527 290147 202561 290175
rect 202589 290147 202623 290175
rect 202651 290147 217797 290175
rect 217825 290147 217859 290175
rect 217887 290147 217921 290175
rect 217949 290147 217983 290175
rect 218011 290147 233157 290175
rect 233185 290147 233219 290175
rect 233247 290147 233281 290175
rect 233309 290147 233343 290175
rect 233371 290147 248517 290175
rect 248545 290147 248579 290175
rect 248607 290147 248641 290175
rect 248669 290147 248703 290175
rect 248731 290147 263877 290175
rect 263905 290147 263939 290175
rect 263967 290147 264001 290175
rect 264029 290147 264063 290175
rect 264091 290147 279237 290175
rect 279265 290147 279299 290175
rect 279327 290147 279361 290175
rect 279389 290147 279423 290175
rect 279451 290147 294597 290175
rect 294625 290147 294659 290175
rect 294687 290147 294721 290175
rect 294749 290147 294783 290175
rect 294811 290147 298248 290175
rect 298276 290147 298310 290175
rect 298338 290147 298372 290175
rect 298400 290147 298434 290175
rect 298462 290147 298990 290175
rect -958 290113 298990 290147
rect -958 290085 -430 290113
rect -402 290085 -368 290113
rect -340 290085 -306 290113
rect -278 290085 -244 290113
rect -216 290085 2757 290113
rect 2785 290085 2819 290113
rect 2847 290085 2881 290113
rect 2909 290085 2943 290113
rect 2971 290085 18117 290113
rect 18145 290085 18179 290113
rect 18207 290085 18241 290113
rect 18269 290085 18303 290113
rect 18331 290085 33477 290113
rect 33505 290085 33539 290113
rect 33567 290085 33601 290113
rect 33629 290085 33663 290113
rect 33691 290085 48837 290113
rect 48865 290085 48899 290113
rect 48927 290085 48961 290113
rect 48989 290085 49023 290113
rect 49051 290085 64197 290113
rect 64225 290085 64259 290113
rect 64287 290085 64321 290113
rect 64349 290085 64383 290113
rect 64411 290085 79557 290113
rect 79585 290085 79619 290113
rect 79647 290085 79681 290113
rect 79709 290085 79743 290113
rect 79771 290085 94917 290113
rect 94945 290085 94979 290113
rect 95007 290085 95041 290113
rect 95069 290085 95103 290113
rect 95131 290085 110277 290113
rect 110305 290085 110339 290113
rect 110367 290085 110401 290113
rect 110429 290085 110463 290113
rect 110491 290085 125637 290113
rect 125665 290085 125699 290113
rect 125727 290085 125761 290113
rect 125789 290085 125823 290113
rect 125851 290085 140997 290113
rect 141025 290085 141059 290113
rect 141087 290085 141121 290113
rect 141149 290085 141183 290113
rect 141211 290085 156357 290113
rect 156385 290085 156419 290113
rect 156447 290085 156481 290113
rect 156509 290085 156543 290113
rect 156571 290085 171717 290113
rect 171745 290085 171779 290113
rect 171807 290085 171841 290113
rect 171869 290085 171903 290113
rect 171931 290085 187077 290113
rect 187105 290085 187139 290113
rect 187167 290085 187201 290113
rect 187229 290085 187263 290113
rect 187291 290085 202437 290113
rect 202465 290085 202499 290113
rect 202527 290085 202561 290113
rect 202589 290085 202623 290113
rect 202651 290085 217797 290113
rect 217825 290085 217859 290113
rect 217887 290085 217921 290113
rect 217949 290085 217983 290113
rect 218011 290085 233157 290113
rect 233185 290085 233219 290113
rect 233247 290085 233281 290113
rect 233309 290085 233343 290113
rect 233371 290085 248517 290113
rect 248545 290085 248579 290113
rect 248607 290085 248641 290113
rect 248669 290085 248703 290113
rect 248731 290085 263877 290113
rect 263905 290085 263939 290113
rect 263967 290085 264001 290113
rect 264029 290085 264063 290113
rect 264091 290085 279237 290113
rect 279265 290085 279299 290113
rect 279327 290085 279361 290113
rect 279389 290085 279423 290113
rect 279451 290085 294597 290113
rect 294625 290085 294659 290113
rect 294687 290085 294721 290113
rect 294749 290085 294783 290113
rect 294811 290085 298248 290113
rect 298276 290085 298310 290113
rect 298338 290085 298372 290113
rect 298400 290085 298434 290113
rect 298462 290085 298990 290113
rect -958 290051 298990 290085
rect -958 290023 -430 290051
rect -402 290023 -368 290051
rect -340 290023 -306 290051
rect -278 290023 -244 290051
rect -216 290023 2757 290051
rect 2785 290023 2819 290051
rect 2847 290023 2881 290051
rect 2909 290023 2943 290051
rect 2971 290023 18117 290051
rect 18145 290023 18179 290051
rect 18207 290023 18241 290051
rect 18269 290023 18303 290051
rect 18331 290023 33477 290051
rect 33505 290023 33539 290051
rect 33567 290023 33601 290051
rect 33629 290023 33663 290051
rect 33691 290023 48837 290051
rect 48865 290023 48899 290051
rect 48927 290023 48961 290051
rect 48989 290023 49023 290051
rect 49051 290023 64197 290051
rect 64225 290023 64259 290051
rect 64287 290023 64321 290051
rect 64349 290023 64383 290051
rect 64411 290023 79557 290051
rect 79585 290023 79619 290051
rect 79647 290023 79681 290051
rect 79709 290023 79743 290051
rect 79771 290023 94917 290051
rect 94945 290023 94979 290051
rect 95007 290023 95041 290051
rect 95069 290023 95103 290051
rect 95131 290023 110277 290051
rect 110305 290023 110339 290051
rect 110367 290023 110401 290051
rect 110429 290023 110463 290051
rect 110491 290023 125637 290051
rect 125665 290023 125699 290051
rect 125727 290023 125761 290051
rect 125789 290023 125823 290051
rect 125851 290023 140997 290051
rect 141025 290023 141059 290051
rect 141087 290023 141121 290051
rect 141149 290023 141183 290051
rect 141211 290023 156357 290051
rect 156385 290023 156419 290051
rect 156447 290023 156481 290051
rect 156509 290023 156543 290051
rect 156571 290023 171717 290051
rect 171745 290023 171779 290051
rect 171807 290023 171841 290051
rect 171869 290023 171903 290051
rect 171931 290023 187077 290051
rect 187105 290023 187139 290051
rect 187167 290023 187201 290051
rect 187229 290023 187263 290051
rect 187291 290023 202437 290051
rect 202465 290023 202499 290051
rect 202527 290023 202561 290051
rect 202589 290023 202623 290051
rect 202651 290023 217797 290051
rect 217825 290023 217859 290051
rect 217887 290023 217921 290051
rect 217949 290023 217983 290051
rect 218011 290023 233157 290051
rect 233185 290023 233219 290051
rect 233247 290023 233281 290051
rect 233309 290023 233343 290051
rect 233371 290023 248517 290051
rect 248545 290023 248579 290051
rect 248607 290023 248641 290051
rect 248669 290023 248703 290051
rect 248731 290023 263877 290051
rect 263905 290023 263939 290051
rect 263967 290023 264001 290051
rect 264029 290023 264063 290051
rect 264091 290023 279237 290051
rect 279265 290023 279299 290051
rect 279327 290023 279361 290051
rect 279389 290023 279423 290051
rect 279451 290023 294597 290051
rect 294625 290023 294659 290051
rect 294687 290023 294721 290051
rect 294749 290023 294783 290051
rect 294811 290023 298248 290051
rect 298276 290023 298310 290051
rect 298338 290023 298372 290051
rect 298400 290023 298434 290051
rect 298462 290023 298990 290051
rect -958 289989 298990 290023
rect -958 289961 -430 289989
rect -402 289961 -368 289989
rect -340 289961 -306 289989
rect -278 289961 -244 289989
rect -216 289961 2757 289989
rect 2785 289961 2819 289989
rect 2847 289961 2881 289989
rect 2909 289961 2943 289989
rect 2971 289961 18117 289989
rect 18145 289961 18179 289989
rect 18207 289961 18241 289989
rect 18269 289961 18303 289989
rect 18331 289961 33477 289989
rect 33505 289961 33539 289989
rect 33567 289961 33601 289989
rect 33629 289961 33663 289989
rect 33691 289961 48837 289989
rect 48865 289961 48899 289989
rect 48927 289961 48961 289989
rect 48989 289961 49023 289989
rect 49051 289961 64197 289989
rect 64225 289961 64259 289989
rect 64287 289961 64321 289989
rect 64349 289961 64383 289989
rect 64411 289961 79557 289989
rect 79585 289961 79619 289989
rect 79647 289961 79681 289989
rect 79709 289961 79743 289989
rect 79771 289961 94917 289989
rect 94945 289961 94979 289989
rect 95007 289961 95041 289989
rect 95069 289961 95103 289989
rect 95131 289961 110277 289989
rect 110305 289961 110339 289989
rect 110367 289961 110401 289989
rect 110429 289961 110463 289989
rect 110491 289961 125637 289989
rect 125665 289961 125699 289989
rect 125727 289961 125761 289989
rect 125789 289961 125823 289989
rect 125851 289961 140997 289989
rect 141025 289961 141059 289989
rect 141087 289961 141121 289989
rect 141149 289961 141183 289989
rect 141211 289961 156357 289989
rect 156385 289961 156419 289989
rect 156447 289961 156481 289989
rect 156509 289961 156543 289989
rect 156571 289961 171717 289989
rect 171745 289961 171779 289989
rect 171807 289961 171841 289989
rect 171869 289961 171903 289989
rect 171931 289961 187077 289989
rect 187105 289961 187139 289989
rect 187167 289961 187201 289989
rect 187229 289961 187263 289989
rect 187291 289961 202437 289989
rect 202465 289961 202499 289989
rect 202527 289961 202561 289989
rect 202589 289961 202623 289989
rect 202651 289961 217797 289989
rect 217825 289961 217859 289989
rect 217887 289961 217921 289989
rect 217949 289961 217983 289989
rect 218011 289961 233157 289989
rect 233185 289961 233219 289989
rect 233247 289961 233281 289989
rect 233309 289961 233343 289989
rect 233371 289961 248517 289989
rect 248545 289961 248579 289989
rect 248607 289961 248641 289989
rect 248669 289961 248703 289989
rect 248731 289961 263877 289989
rect 263905 289961 263939 289989
rect 263967 289961 264001 289989
rect 264029 289961 264063 289989
rect 264091 289961 279237 289989
rect 279265 289961 279299 289989
rect 279327 289961 279361 289989
rect 279389 289961 279423 289989
rect 279451 289961 294597 289989
rect 294625 289961 294659 289989
rect 294687 289961 294721 289989
rect 294749 289961 294783 289989
rect 294811 289961 298248 289989
rect 298276 289961 298310 289989
rect 298338 289961 298372 289989
rect 298400 289961 298434 289989
rect 298462 289961 298990 289989
rect -958 289913 298990 289961
rect -958 284175 298990 284223
rect -958 284147 -910 284175
rect -882 284147 -848 284175
rect -820 284147 -786 284175
rect -758 284147 -724 284175
rect -696 284147 4617 284175
rect 4645 284147 4679 284175
rect 4707 284147 4741 284175
rect 4769 284147 4803 284175
rect 4831 284147 19977 284175
rect 20005 284147 20039 284175
rect 20067 284147 20101 284175
rect 20129 284147 20163 284175
rect 20191 284147 35337 284175
rect 35365 284147 35399 284175
rect 35427 284147 35461 284175
rect 35489 284147 35523 284175
rect 35551 284147 50697 284175
rect 50725 284147 50759 284175
rect 50787 284147 50821 284175
rect 50849 284147 50883 284175
rect 50911 284147 66057 284175
rect 66085 284147 66119 284175
rect 66147 284147 66181 284175
rect 66209 284147 66243 284175
rect 66271 284147 81417 284175
rect 81445 284147 81479 284175
rect 81507 284147 81541 284175
rect 81569 284147 81603 284175
rect 81631 284147 96777 284175
rect 96805 284147 96839 284175
rect 96867 284147 96901 284175
rect 96929 284147 96963 284175
rect 96991 284147 112137 284175
rect 112165 284147 112199 284175
rect 112227 284147 112261 284175
rect 112289 284147 112323 284175
rect 112351 284147 127497 284175
rect 127525 284147 127559 284175
rect 127587 284147 127621 284175
rect 127649 284147 127683 284175
rect 127711 284147 142857 284175
rect 142885 284147 142919 284175
rect 142947 284147 142981 284175
rect 143009 284147 143043 284175
rect 143071 284147 158217 284175
rect 158245 284147 158279 284175
rect 158307 284147 158341 284175
rect 158369 284147 158403 284175
rect 158431 284147 173577 284175
rect 173605 284147 173639 284175
rect 173667 284147 173701 284175
rect 173729 284147 173763 284175
rect 173791 284147 188937 284175
rect 188965 284147 188999 284175
rect 189027 284147 189061 284175
rect 189089 284147 189123 284175
rect 189151 284147 204297 284175
rect 204325 284147 204359 284175
rect 204387 284147 204421 284175
rect 204449 284147 204483 284175
rect 204511 284147 219657 284175
rect 219685 284147 219719 284175
rect 219747 284147 219781 284175
rect 219809 284147 219843 284175
rect 219871 284147 235017 284175
rect 235045 284147 235079 284175
rect 235107 284147 235141 284175
rect 235169 284147 235203 284175
rect 235231 284147 250377 284175
rect 250405 284147 250439 284175
rect 250467 284147 250501 284175
rect 250529 284147 250563 284175
rect 250591 284147 265737 284175
rect 265765 284147 265799 284175
rect 265827 284147 265861 284175
rect 265889 284147 265923 284175
rect 265951 284147 281097 284175
rect 281125 284147 281159 284175
rect 281187 284147 281221 284175
rect 281249 284147 281283 284175
rect 281311 284147 296457 284175
rect 296485 284147 296519 284175
rect 296547 284147 296581 284175
rect 296609 284147 296643 284175
rect 296671 284147 298728 284175
rect 298756 284147 298790 284175
rect 298818 284147 298852 284175
rect 298880 284147 298914 284175
rect 298942 284147 298990 284175
rect -958 284113 298990 284147
rect -958 284085 -910 284113
rect -882 284085 -848 284113
rect -820 284085 -786 284113
rect -758 284085 -724 284113
rect -696 284085 4617 284113
rect 4645 284085 4679 284113
rect 4707 284085 4741 284113
rect 4769 284085 4803 284113
rect 4831 284085 19977 284113
rect 20005 284085 20039 284113
rect 20067 284085 20101 284113
rect 20129 284085 20163 284113
rect 20191 284085 35337 284113
rect 35365 284085 35399 284113
rect 35427 284085 35461 284113
rect 35489 284085 35523 284113
rect 35551 284085 50697 284113
rect 50725 284085 50759 284113
rect 50787 284085 50821 284113
rect 50849 284085 50883 284113
rect 50911 284085 66057 284113
rect 66085 284085 66119 284113
rect 66147 284085 66181 284113
rect 66209 284085 66243 284113
rect 66271 284085 81417 284113
rect 81445 284085 81479 284113
rect 81507 284085 81541 284113
rect 81569 284085 81603 284113
rect 81631 284085 96777 284113
rect 96805 284085 96839 284113
rect 96867 284085 96901 284113
rect 96929 284085 96963 284113
rect 96991 284085 112137 284113
rect 112165 284085 112199 284113
rect 112227 284085 112261 284113
rect 112289 284085 112323 284113
rect 112351 284085 127497 284113
rect 127525 284085 127559 284113
rect 127587 284085 127621 284113
rect 127649 284085 127683 284113
rect 127711 284085 142857 284113
rect 142885 284085 142919 284113
rect 142947 284085 142981 284113
rect 143009 284085 143043 284113
rect 143071 284085 158217 284113
rect 158245 284085 158279 284113
rect 158307 284085 158341 284113
rect 158369 284085 158403 284113
rect 158431 284085 173577 284113
rect 173605 284085 173639 284113
rect 173667 284085 173701 284113
rect 173729 284085 173763 284113
rect 173791 284085 188937 284113
rect 188965 284085 188999 284113
rect 189027 284085 189061 284113
rect 189089 284085 189123 284113
rect 189151 284085 204297 284113
rect 204325 284085 204359 284113
rect 204387 284085 204421 284113
rect 204449 284085 204483 284113
rect 204511 284085 219657 284113
rect 219685 284085 219719 284113
rect 219747 284085 219781 284113
rect 219809 284085 219843 284113
rect 219871 284085 235017 284113
rect 235045 284085 235079 284113
rect 235107 284085 235141 284113
rect 235169 284085 235203 284113
rect 235231 284085 250377 284113
rect 250405 284085 250439 284113
rect 250467 284085 250501 284113
rect 250529 284085 250563 284113
rect 250591 284085 265737 284113
rect 265765 284085 265799 284113
rect 265827 284085 265861 284113
rect 265889 284085 265923 284113
rect 265951 284085 281097 284113
rect 281125 284085 281159 284113
rect 281187 284085 281221 284113
rect 281249 284085 281283 284113
rect 281311 284085 296457 284113
rect 296485 284085 296519 284113
rect 296547 284085 296581 284113
rect 296609 284085 296643 284113
rect 296671 284085 298728 284113
rect 298756 284085 298790 284113
rect 298818 284085 298852 284113
rect 298880 284085 298914 284113
rect 298942 284085 298990 284113
rect -958 284051 298990 284085
rect -958 284023 -910 284051
rect -882 284023 -848 284051
rect -820 284023 -786 284051
rect -758 284023 -724 284051
rect -696 284023 4617 284051
rect 4645 284023 4679 284051
rect 4707 284023 4741 284051
rect 4769 284023 4803 284051
rect 4831 284023 19977 284051
rect 20005 284023 20039 284051
rect 20067 284023 20101 284051
rect 20129 284023 20163 284051
rect 20191 284023 35337 284051
rect 35365 284023 35399 284051
rect 35427 284023 35461 284051
rect 35489 284023 35523 284051
rect 35551 284023 50697 284051
rect 50725 284023 50759 284051
rect 50787 284023 50821 284051
rect 50849 284023 50883 284051
rect 50911 284023 66057 284051
rect 66085 284023 66119 284051
rect 66147 284023 66181 284051
rect 66209 284023 66243 284051
rect 66271 284023 81417 284051
rect 81445 284023 81479 284051
rect 81507 284023 81541 284051
rect 81569 284023 81603 284051
rect 81631 284023 96777 284051
rect 96805 284023 96839 284051
rect 96867 284023 96901 284051
rect 96929 284023 96963 284051
rect 96991 284023 112137 284051
rect 112165 284023 112199 284051
rect 112227 284023 112261 284051
rect 112289 284023 112323 284051
rect 112351 284023 127497 284051
rect 127525 284023 127559 284051
rect 127587 284023 127621 284051
rect 127649 284023 127683 284051
rect 127711 284023 142857 284051
rect 142885 284023 142919 284051
rect 142947 284023 142981 284051
rect 143009 284023 143043 284051
rect 143071 284023 158217 284051
rect 158245 284023 158279 284051
rect 158307 284023 158341 284051
rect 158369 284023 158403 284051
rect 158431 284023 173577 284051
rect 173605 284023 173639 284051
rect 173667 284023 173701 284051
rect 173729 284023 173763 284051
rect 173791 284023 188937 284051
rect 188965 284023 188999 284051
rect 189027 284023 189061 284051
rect 189089 284023 189123 284051
rect 189151 284023 204297 284051
rect 204325 284023 204359 284051
rect 204387 284023 204421 284051
rect 204449 284023 204483 284051
rect 204511 284023 219657 284051
rect 219685 284023 219719 284051
rect 219747 284023 219781 284051
rect 219809 284023 219843 284051
rect 219871 284023 235017 284051
rect 235045 284023 235079 284051
rect 235107 284023 235141 284051
rect 235169 284023 235203 284051
rect 235231 284023 250377 284051
rect 250405 284023 250439 284051
rect 250467 284023 250501 284051
rect 250529 284023 250563 284051
rect 250591 284023 265737 284051
rect 265765 284023 265799 284051
rect 265827 284023 265861 284051
rect 265889 284023 265923 284051
rect 265951 284023 281097 284051
rect 281125 284023 281159 284051
rect 281187 284023 281221 284051
rect 281249 284023 281283 284051
rect 281311 284023 296457 284051
rect 296485 284023 296519 284051
rect 296547 284023 296581 284051
rect 296609 284023 296643 284051
rect 296671 284023 298728 284051
rect 298756 284023 298790 284051
rect 298818 284023 298852 284051
rect 298880 284023 298914 284051
rect 298942 284023 298990 284051
rect -958 283989 298990 284023
rect -958 283961 -910 283989
rect -882 283961 -848 283989
rect -820 283961 -786 283989
rect -758 283961 -724 283989
rect -696 283961 4617 283989
rect 4645 283961 4679 283989
rect 4707 283961 4741 283989
rect 4769 283961 4803 283989
rect 4831 283961 19977 283989
rect 20005 283961 20039 283989
rect 20067 283961 20101 283989
rect 20129 283961 20163 283989
rect 20191 283961 35337 283989
rect 35365 283961 35399 283989
rect 35427 283961 35461 283989
rect 35489 283961 35523 283989
rect 35551 283961 50697 283989
rect 50725 283961 50759 283989
rect 50787 283961 50821 283989
rect 50849 283961 50883 283989
rect 50911 283961 66057 283989
rect 66085 283961 66119 283989
rect 66147 283961 66181 283989
rect 66209 283961 66243 283989
rect 66271 283961 81417 283989
rect 81445 283961 81479 283989
rect 81507 283961 81541 283989
rect 81569 283961 81603 283989
rect 81631 283961 96777 283989
rect 96805 283961 96839 283989
rect 96867 283961 96901 283989
rect 96929 283961 96963 283989
rect 96991 283961 112137 283989
rect 112165 283961 112199 283989
rect 112227 283961 112261 283989
rect 112289 283961 112323 283989
rect 112351 283961 127497 283989
rect 127525 283961 127559 283989
rect 127587 283961 127621 283989
rect 127649 283961 127683 283989
rect 127711 283961 142857 283989
rect 142885 283961 142919 283989
rect 142947 283961 142981 283989
rect 143009 283961 143043 283989
rect 143071 283961 158217 283989
rect 158245 283961 158279 283989
rect 158307 283961 158341 283989
rect 158369 283961 158403 283989
rect 158431 283961 173577 283989
rect 173605 283961 173639 283989
rect 173667 283961 173701 283989
rect 173729 283961 173763 283989
rect 173791 283961 188937 283989
rect 188965 283961 188999 283989
rect 189027 283961 189061 283989
rect 189089 283961 189123 283989
rect 189151 283961 204297 283989
rect 204325 283961 204359 283989
rect 204387 283961 204421 283989
rect 204449 283961 204483 283989
rect 204511 283961 219657 283989
rect 219685 283961 219719 283989
rect 219747 283961 219781 283989
rect 219809 283961 219843 283989
rect 219871 283961 235017 283989
rect 235045 283961 235079 283989
rect 235107 283961 235141 283989
rect 235169 283961 235203 283989
rect 235231 283961 250377 283989
rect 250405 283961 250439 283989
rect 250467 283961 250501 283989
rect 250529 283961 250563 283989
rect 250591 283961 265737 283989
rect 265765 283961 265799 283989
rect 265827 283961 265861 283989
rect 265889 283961 265923 283989
rect 265951 283961 281097 283989
rect 281125 283961 281159 283989
rect 281187 283961 281221 283989
rect 281249 283961 281283 283989
rect 281311 283961 296457 283989
rect 296485 283961 296519 283989
rect 296547 283961 296581 283989
rect 296609 283961 296643 283989
rect 296671 283961 298728 283989
rect 298756 283961 298790 283989
rect 298818 283961 298852 283989
rect 298880 283961 298914 283989
rect 298942 283961 298990 283989
rect -958 283913 298990 283961
rect -958 281175 298990 281223
rect -958 281147 -430 281175
rect -402 281147 -368 281175
rect -340 281147 -306 281175
rect -278 281147 -244 281175
rect -216 281147 2757 281175
rect 2785 281147 2819 281175
rect 2847 281147 2881 281175
rect 2909 281147 2943 281175
rect 2971 281147 18117 281175
rect 18145 281147 18179 281175
rect 18207 281147 18241 281175
rect 18269 281147 18303 281175
rect 18331 281147 33477 281175
rect 33505 281147 33539 281175
rect 33567 281147 33601 281175
rect 33629 281147 33663 281175
rect 33691 281147 48837 281175
rect 48865 281147 48899 281175
rect 48927 281147 48961 281175
rect 48989 281147 49023 281175
rect 49051 281147 64197 281175
rect 64225 281147 64259 281175
rect 64287 281147 64321 281175
rect 64349 281147 64383 281175
rect 64411 281147 79557 281175
rect 79585 281147 79619 281175
rect 79647 281147 79681 281175
rect 79709 281147 79743 281175
rect 79771 281147 94917 281175
rect 94945 281147 94979 281175
rect 95007 281147 95041 281175
rect 95069 281147 95103 281175
rect 95131 281147 110277 281175
rect 110305 281147 110339 281175
rect 110367 281147 110401 281175
rect 110429 281147 110463 281175
rect 110491 281147 125637 281175
rect 125665 281147 125699 281175
rect 125727 281147 125761 281175
rect 125789 281147 125823 281175
rect 125851 281147 140997 281175
rect 141025 281147 141059 281175
rect 141087 281147 141121 281175
rect 141149 281147 141183 281175
rect 141211 281147 156357 281175
rect 156385 281147 156419 281175
rect 156447 281147 156481 281175
rect 156509 281147 156543 281175
rect 156571 281147 171717 281175
rect 171745 281147 171779 281175
rect 171807 281147 171841 281175
rect 171869 281147 171903 281175
rect 171931 281147 187077 281175
rect 187105 281147 187139 281175
rect 187167 281147 187201 281175
rect 187229 281147 187263 281175
rect 187291 281147 202437 281175
rect 202465 281147 202499 281175
rect 202527 281147 202561 281175
rect 202589 281147 202623 281175
rect 202651 281147 217797 281175
rect 217825 281147 217859 281175
rect 217887 281147 217921 281175
rect 217949 281147 217983 281175
rect 218011 281147 233157 281175
rect 233185 281147 233219 281175
rect 233247 281147 233281 281175
rect 233309 281147 233343 281175
rect 233371 281147 248517 281175
rect 248545 281147 248579 281175
rect 248607 281147 248641 281175
rect 248669 281147 248703 281175
rect 248731 281147 263877 281175
rect 263905 281147 263939 281175
rect 263967 281147 264001 281175
rect 264029 281147 264063 281175
rect 264091 281147 279237 281175
rect 279265 281147 279299 281175
rect 279327 281147 279361 281175
rect 279389 281147 279423 281175
rect 279451 281147 294597 281175
rect 294625 281147 294659 281175
rect 294687 281147 294721 281175
rect 294749 281147 294783 281175
rect 294811 281147 298248 281175
rect 298276 281147 298310 281175
rect 298338 281147 298372 281175
rect 298400 281147 298434 281175
rect 298462 281147 298990 281175
rect -958 281113 298990 281147
rect -958 281085 -430 281113
rect -402 281085 -368 281113
rect -340 281085 -306 281113
rect -278 281085 -244 281113
rect -216 281085 2757 281113
rect 2785 281085 2819 281113
rect 2847 281085 2881 281113
rect 2909 281085 2943 281113
rect 2971 281085 18117 281113
rect 18145 281085 18179 281113
rect 18207 281085 18241 281113
rect 18269 281085 18303 281113
rect 18331 281085 33477 281113
rect 33505 281085 33539 281113
rect 33567 281085 33601 281113
rect 33629 281085 33663 281113
rect 33691 281085 48837 281113
rect 48865 281085 48899 281113
rect 48927 281085 48961 281113
rect 48989 281085 49023 281113
rect 49051 281085 64197 281113
rect 64225 281085 64259 281113
rect 64287 281085 64321 281113
rect 64349 281085 64383 281113
rect 64411 281085 79557 281113
rect 79585 281085 79619 281113
rect 79647 281085 79681 281113
rect 79709 281085 79743 281113
rect 79771 281085 94917 281113
rect 94945 281085 94979 281113
rect 95007 281085 95041 281113
rect 95069 281085 95103 281113
rect 95131 281085 110277 281113
rect 110305 281085 110339 281113
rect 110367 281085 110401 281113
rect 110429 281085 110463 281113
rect 110491 281085 125637 281113
rect 125665 281085 125699 281113
rect 125727 281085 125761 281113
rect 125789 281085 125823 281113
rect 125851 281085 140997 281113
rect 141025 281085 141059 281113
rect 141087 281085 141121 281113
rect 141149 281085 141183 281113
rect 141211 281085 156357 281113
rect 156385 281085 156419 281113
rect 156447 281085 156481 281113
rect 156509 281085 156543 281113
rect 156571 281085 171717 281113
rect 171745 281085 171779 281113
rect 171807 281085 171841 281113
rect 171869 281085 171903 281113
rect 171931 281085 187077 281113
rect 187105 281085 187139 281113
rect 187167 281085 187201 281113
rect 187229 281085 187263 281113
rect 187291 281085 202437 281113
rect 202465 281085 202499 281113
rect 202527 281085 202561 281113
rect 202589 281085 202623 281113
rect 202651 281085 217797 281113
rect 217825 281085 217859 281113
rect 217887 281085 217921 281113
rect 217949 281085 217983 281113
rect 218011 281085 233157 281113
rect 233185 281085 233219 281113
rect 233247 281085 233281 281113
rect 233309 281085 233343 281113
rect 233371 281085 248517 281113
rect 248545 281085 248579 281113
rect 248607 281085 248641 281113
rect 248669 281085 248703 281113
rect 248731 281085 263877 281113
rect 263905 281085 263939 281113
rect 263967 281085 264001 281113
rect 264029 281085 264063 281113
rect 264091 281085 279237 281113
rect 279265 281085 279299 281113
rect 279327 281085 279361 281113
rect 279389 281085 279423 281113
rect 279451 281085 294597 281113
rect 294625 281085 294659 281113
rect 294687 281085 294721 281113
rect 294749 281085 294783 281113
rect 294811 281085 298248 281113
rect 298276 281085 298310 281113
rect 298338 281085 298372 281113
rect 298400 281085 298434 281113
rect 298462 281085 298990 281113
rect -958 281051 298990 281085
rect -958 281023 -430 281051
rect -402 281023 -368 281051
rect -340 281023 -306 281051
rect -278 281023 -244 281051
rect -216 281023 2757 281051
rect 2785 281023 2819 281051
rect 2847 281023 2881 281051
rect 2909 281023 2943 281051
rect 2971 281023 18117 281051
rect 18145 281023 18179 281051
rect 18207 281023 18241 281051
rect 18269 281023 18303 281051
rect 18331 281023 33477 281051
rect 33505 281023 33539 281051
rect 33567 281023 33601 281051
rect 33629 281023 33663 281051
rect 33691 281023 48837 281051
rect 48865 281023 48899 281051
rect 48927 281023 48961 281051
rect 48989 281023 49023 281051
rect 49051 281023 64197 281051
rect 64225 281023 64259 281051
rect 64287 281023 64321 281051
rect 64349 281023 64383 281051
rect 64411 281023 79557 281051
rect 79585 281023 79619 281051
rect 79647 281023 79681 281051
rect 79709 281023 79743 281051
rect 79771 281023 94917 281051
rect 94945 281023 94979 281051
rect 95007 281023 95041 281051
rect 95069 281023 95103 281051
rect 95131 281023 110277 281051
rect 110305 281023 110339 281051
rect 110367 281023 110401 281051
rect 110429 281023 110463 281051
rect 110491 281023 125637 281051
rect 125665 281023 125699 281051
rect 125727 281023 125761 281051
rect 125789 281023 125823 281051
rect 125851 281023 140997 281051
rect 141025 281023 141059 281051
rect 141087 281023 141121 281051
rect 141149 281023 141183 281051
rect 141211 281023 156357 281051
rect 156385 281023 156419 281051
rect 156447 281023 156481 281051
rect 156509 281023 156543 281051
rect 156571 281023 171717 281051
rect 171745 281023 171779 281051
rect 171807 281023 171841 281051
rect 171869 281023 171903 281051
rect 171931 281023 187077 281051
rect 187105 281023 187139 281051
rect 187167 281023 187201 281051
rect 187229 281023 187263 281051
rect 187291 281023 202437 281051
rect 202465 281023 202499 281051
rect 202527 281023 202561 281051
rect 202589 281023 202623 281051
rect 202651 281023 217797 281051
rect 217825 281023 217859 281051
rect 217887 281023 217921 281051
rect 217949 281023 217983 281051
rect 218011 281023 233157 281051
rect 233185 281023 233219 281051
rect 233247 281023 233281 281051
rect 233309 281023 233343 281051
rect 233371 281023 248517 281051
rect 248545 281023 248579 281051
rect 248607 281023 248641 281051
rect 248669 281023 248703 281051
rect 248731 281023 263877 281051
rect 263905 281023 263939 281051
rect 263967 281023 264001 281051
rect 264029 281023 264063 281051
rect 264091 281023 279237 281051
rect 279265 281023 279299 281051
rect 279327 281023 279361 281051
rect 279389 281023 279423 281051
rect 279451 281023 294597 281051
rect 294625 281023 294659 281051
rect 294687 281023 294721 281051
rect 294749 281023 294783 281051
rect 294811 281023 298248 281051
rect 298276 281023 298310 281051
rect 298338 281023 298372 281051
rect 298400 281023 298434 281051
rect 298462 281023 298990 281051
rect -958 280989 298990 281023
rect -958 280961 -430 280989
rect -402 280961 -368 280989
rect -340 280961 -306 280989
rect -278 280961 -244 280989
rect -216 280961 2757 280989
rect 2785 280961 2819 280989
rect 2847 280961 2881 280989
rect 2909 280961 2943 280989
rect 2971 280961 18117 280989
rect 18145 280961 18179 280989
rect 18207 280961 18241 280989
rect 18269 280961 18303 280989
rect 18331 280961 33477 280989
rect 33505 280961 33539 280989
rect 33567 280961 33601 280989
rect 33629 280961 33663 280989
rect 33691 280961 48837 280989
rect 48865 280961 48899 280989
rect 48927 280961 48961 280989
rect 48989 280961 49023 280989
rect 49051 280961 64197 280989
rect 64225 280961 64259 280989
rect 64287 280961 64321 280989
rect 64349 280961 64383 280989
rect 64411 280961 79557 280989
rect 79585 280961 79619 280989
rect 79647 280961 79681 280989
rect 79709 280961 79743 280989
rect 79771 280961 94917 280989
rect 94945 280961 94979 280989
rect 95007 280961 95041 280989
rect 95069 280961 95103 280989
rect 95131 280961 110277 280989
rect 110305 280961 110339 280989
rect 110367 280961 110401 280989
rect 110429 280961 110463 280989
rect 110491 280961 125637 280989
rect 125665 280961 125699 280989
rect 125727 280961 125761 280989
rect 125789 280961 125823 280989
rect 125851 280961 140997 280989
rect 141025 280961 141059 280989
rect 141087 280961 141121 280989
rect 141149 280961 141183 280989
rect 141211 280961 156357 280989
rect 156385 280961 156419 280989
rect 156447 280961 156481 280989
rect 156509 280961 156543 280989
rect 156571 280961 171717 280989
rect 171745 280961 171779 280989
rect 171807 280961 171841 280989
rect 171869 280961 171903 280989
rect 171931 280961 187077 280989
rect 187105 280961 187139 280989
rect 187167 280961 187201 280989
rect 187229 280961 187263 280989
rect 187291 280961 202437 280989
rect 202465 280961 202499 280989
rect 202527 280961 202561 280989
rect 202589 280961 202623 280989
rect 202651 280961 217797 280989
rect 217825 280961 217859 280989
rect 217887 280961 217921 280989
rect 217949 280961 217983 280989
rect 218011 280961 233157 280989
rect 233185 280961 233219 280989
rect 233247 280961 233281 280989
rect 233309 280961 233343 280989
rect 233371 280961 248517 280989
rect 248545 280961 248579 280989
rect 248607 280961 248641 280989
rect 248669 280961 248703 280989
rect 248731 280961 263877 280989
rect 263905 280961 263939 280989
rect 263967 280961 264001 280989
rect 264029 280961 264063 280989
rect 264091 280961 279237 280989
rect 279265 280961 279299 280989
rect 279327 280961 279361 280989
rect 279389 280961 279423 280989
rect 279451 280961 294597 280989
rect 294625 280961 294659 280989
rect 294687 280961 294721 280989
rect 294749 280961 294783 280989
rect 294811 280961 298248 280989
rect 298276 280961 298310 280989
rect 298338 280961 298372 280989
rect 298400 280961 298434 280989
rect 298462 280961 298990 280989
rect -958 280913 298990 280961
rect -958 275175 298990 275223
rect -958 275147 -910 275175
rect -882 275147 -848 275175
rect -820 275147 -786 275175
rect -758 275147 -724 275175
rect -696 275147 4617 275175
rect 4645 275147 4679 275175
rect 4707 275147 4741 275175
rect 4769 275147 4803 275175
rect 4831 275147 19977 275175
rect 20005 275147 20039 275175
rect 20067 275147 20101 275175
rect 20129 275147 20163 275175
rect 20191 275147 35337 275175
rect 35365 275147 35399 275175
rect 35427 275147 35461 275175
rect 35489 275147 35523 275175
rect 35551 275147 50697 275175
rect 50725 275147 50759 275175
rect 50787 275147 50821 275175
rect 50849 275147 50883 275175
rect 50911 275147 66057 275175
rect 66085 275147 66119 275175
rect 66147 275147 66181 275175
rect 66209 275147 66243 275175
rect 66271 275147 81417 275175
rect 81445 275147 81479 275175
rect 81507 275147 81541 275175
rect 81569 275147 81603 275175
rect 81631 275147 96777 275175
rect 96805 275147 96839 275175
rect 96867 275147 96901 275175
rect 96929 275147 96963 275175
rect 96991 275147 112137 275175
rect 112165 275147 112199 275175
rect 112227 275147 112261 275175
rect 112289 275147 112323 275175
rect 112351 275147 127497 275175
rect 127525 275147 127559 275175
rect 127587 275147 127621 275175
rect 127649 275147 127683 275175
rect 127711 275147 142857 275175
rect 142885 275147 142919 275175
rect 142947 275147 142981 275175
rect 143009 275147 143043 275175
rect 143071 275147 158217 275175
rect 158245 275147 158279 275175
rect 158307 275147 158341 275175
rect 158369 275147 158403 275175
rect 158431 275147 173577 275175
rect 173605 275147 173639 275175
rect 173667 275147 173701 275175
rect 173729 275147 173763 275175
rect 173791 275147 188937 275175
rect 188965 275147 188999 275175
rect 189027 275147 189061 275175
rect 189089 275147 189123 275175
rect 189151 275147 204297 275175
rect 204325 275147 204359 275175
rect 204387 275147 204421 275175
rect 204449 275147 204483 275175
rect 204511 275147 219657 275175
rect 219685 275147 219719 275175
rect 219747 275147 219781 275175
rect 219809 275147 219843 275175
rect 219871 275147 235017 275175
rect 235045 275147 235079 275175
rect 235107 275147 235141 275175
rect 235169 275147 235203 275175
rect 235231 275147 250377 275175
rect 250405 275147 250439 275175
rect 250467 275147 250501 275175
rect 250529 275147 250563 275175
rect 250591 275147 265737 275175
rect 265765 275147 265799 275175
rect 265827 275147 265861 275175
rect 265889 275147 265923 275175
rect 265951 275147 281097 275175
rect 281125 275147 281159 275175
rect 281187 275147 281221 275175
rect 281249 275147 281283 275175
rect 281311 275147 296457 275175
rect 296485 275147 296519 275175
rect 296547 275147 296581 275175
rect 296609 275147 296643 275175
rect 296671 275147 298728 275175
rect 298756 275147 298790 275175
rect 298818 275147 298852 275175
rect 298880 275147 298914 275175
rect 298942 275147 298990 275175
rect -958 275113 298990 275147
rect -958 275085 -910 275113
rect -882 275085 -848 275113
rect -820 275085 -786 275113
rect -758 275085 -724 275113
rect -696 275085 4617 275113
rect 4645 275085 4679 275113
rect 4707 275085 4741 275113
rect 4769 275085 4803 275113
rect 4831 275085 19977 275113
rect 20005 275085 20039 275113
rect 20067 275085 20101 275113
rect 20129 275085 20163 275113
rect 20191 275085 35337 275113
rect 35365 275085 35399 275113
rect 35427 275085 35461 275113
rect 35489 275085 35523 275113
rect 35551 275085 50697 275113
rect 50725 275085 50759 275113
rect 50787 275085 50821 275113
rect 50849 275085 50883 275113
rect 50911 275085 66057 275113
rect 66085 275085 66119 275113
rect 66147 275085 66181 275113
rect 66209 275085 66243 275113
rect 66271 275085 81417 275113
rect 81445 275085 81479 275113
rect 81507 275085 81541 275113
rect 81569 275085 81603 275113
rect 81631 275085 96777 275113
rect 96805 275085 96839 275113
rect 96867 275085 96901 275113
rect 96929 275085 96963 275113
rect 96991 275085 112137 275113
rect 112165 275085 112199 275113
rect 112227 275085 112261 275113
rect 112289 275085 112323 275113
rect 112351 275085 127497 275113
rect 127525 275085 127559 275113
rect 127587 275085 127621 275113
rect 127649 275085 127683 275113
rect 127711 275085 142857 275113
rect 142885 275085 142919 275113
rect 142947 275085 142981 275113
rect 143009 275085 143043 275113
rect 143071 275085 158217 275113
rect 158245 275085 158279 275113
rect 158307 275085 158341 275113
rect 158369 275085 158403 275113
rect 158431 275085 173577 275113
rect 173605 275085 173639 275113
rect 173667 275085 173701 275113
rect 173729 275085 173763 275113
rect 173791 275085 188937 275113
rect 188965 275085 188999 275113
rect 189027 275085 189061 275113
rect 189089 275085 189123 275113
rect 189151 275085 204297 275113
rect 204325 275085 204359 275113
rect 204387 275085 204421 275113
rect 204449 275085 204483 275113
rect 204511 275085 219657 275113
rect 219685 275085 219719 275113
rect 219747 275085 219781 275113
rect 219809 275085 219843 275113
rect 219871 275085 235017 275113
rect 235045 275085 235079 275113
rect 235107 275085 235141 275113
rect 235169 275085 235203 275113
rect 235231 275085 250377 275113
rect 250405 275085 250439 275113
rect 250467 275085 250501 275113
rect 250529 275085 250563 275113
rect 250591 275085 265737 275113
rect 265765 275085 265799 275113
rect 265827 275085 265861 275113
rect 265889 275085 265923 275113
rect 265951 275085 281097 275113
rect 281125 275085 281159 275113
rect 281187 275085 281221 275113
rect 281249 275085 281283 275113
rect 281311 275085 296457 275113
rect 296485 275085 296519 275113
rect 296547 275085 296581 275113
rect 296609 275085 296643 275113
rect 296671 275085 298728 275113
rect 298756 275085 298790 275113
rect 298818 275085 298852 275113
rect 298880 275085 298914 275113
rect 298942 275085 298990 275113
rect -958 275051 298990 275085
rect -958 275023 -910 275051
rect -882 275023 -848 275051
rect -820 275023 -786 275051
rect -758 275023 -724 275051
rect -696 275023 4617 275051
rect 4645 275023 4679 275051
rect 4707 275023 4741 275051
rect 4769 275023 4803 275051
rect 4831 275023 19977 275051
rect 20005 275023 20039 275051
rect 20067 275023 20101 275051
rect 20129 275023 20163 275051
rect 20191 275023 35337 275051
rect 35365 275023 35399 275051
rect 35427 275023 35461 275051
rect 35489 275023 35523 275051
rect 35551 275023 50697 275051
rect 50725 275023 50759 275051
rect 50787 275023 50821 275051
rect 50849 275023 50883 275051
rect 50911 275023 66057 275051
rect 66085 275023 66119 275051
rect 66147 275023 66181 275051
rect 66209 275023 66243 275051
rect 66271 275023 81417 275051
rect 81445 275023 81479 275051
rect 81507 275023 81541 275051
rect 81569 275023 81603 275051
rect 81631 275023 96777 275051
rect 96805 275023 96839 275051
rect 96867 275023 96901 275051
rect 96929 275023 96963 275051
rect 96991 275023 112137 275051
rect 112165 275023 112199 275051
rect 112227 275023 112261 275051
rect 112289 275023 112323 275051
rect 112351 275023 127497 275051
rect 127525 275023 127559 275051
rect 127587 275023 127621 275051
rect 127649 275023 127683 275051
rect 127711 275023 142857 275051
rect 142885 275023 142919 275051
rect 142947 275023 142981 275051
rect 143009 275023 143043 275051
rect 143071 275023 158217 275051
rect 158245 275023 158279 275051
rect 158307 275023 158341 275051
rect 158369 275023 158403 275051
rect 158431 275023 173577 275051
rect 173605 275023 173639 275051
rect 173667 275023 173701 275051
rect 173729 275023 173763 275051
rect 173791 275023 188937 275051
rect 188965 275023 188999 275051
rect 189027 275023 189061 275051
rect 189089 275023 189123 275051
rect 189151 275023 204297 275051
rect 204325 275023 204359 275051
rect 204387 275023 204421 275051
rect 204449 275023 204483 275051
rect 204511 275023 219657 275051
rect 219685 275023 219719 275051
rect 219747 275023 219781 275051
rect 219809 275023 219843 275051
rect 219871 275023 235017 275051
rect 235045 275023 235079 275051
rect 235107 275023 235141 275051
rect 235169 275023 235203 275051
rect 235231 275023 250377 275051
rect 250405 275023 250439 275051
rect 250467 275023 250501 275051
rect 250529 275023 250563 275051
rect 250591 275023 265737 275051
rect 265765 275023 265799 275051
rect 265827 275023 265861 275051
rect 265889 275023 265923 275051
rect 265951 275023 281097 275051
rect 281125 275023 281159 275051
rect 281187 275023 281221 275051
rect 281249 275023 281283 275051
rect 281311 275023 296457 275051
rect 296485 275023 296519 275051
rect 296547 275023 296581 275051
rect 296609 275023 296643 275051
rect 296671 275023 298728 275051
rect 298756 275023 298790 275051
rect 298818 275023 298852 275051
rect 298880 275023 298914 275051
rect 298942 275023 298990 275051
rect -958 274989 298990 275023
rect -958 274961 -910 274989
rect -882 274961 -848 274989
rect -820 274961 -786 274989
rect -758 274961 -724 274989
rect -696 274961 4617 274989
rect 4645 274961 4679 274989
rect 4707 274961 4741 274989
rect 4769 274961 4803 274989
rect 4831 274961 19977 274989
rect 20005 274961 20039 274989
rect 20067 274961 20101 274989
rect 20129 274961 20163 274989
rect 20191 274961 35337 274989
rect 35365 274961 35399 274989
rect 35427 274961 35461 274989
rect 35489 274961 35523 274989
rect 35551 274961 50697 274989
rect 50725 274961 50759 274989
rect 50787 274961 50821 274989
rect 50849 274961 50883 274989
rect 50911 274961 66057 274989
rect 66085 274961 66119 274989
rect 66147 274961 66181 274989
rect 66209 274961 66243 274989
rect 66271 274961 81417 274989
rect 81445 274961 81479 274989
rect 81507 274961 81541 274989
rect 81569 274961 81603 274989
rect 81631 274961 96777 274989
rect 96805 274961 96839 274989
rect 96867 274961 96901 274989
rect 96929 274961 96963 274989
rect 96991 274961 112137 274989
rect 112165 274961 112199 274989
rect 112227 274961 112261 274989
rect 112289 274961 112323 274989
rect 112351 274961 127497 274989
rect 127525 274961 127559 274989
rect 127587 274961 127621 274989
rect 127649 274961 127683 274989
rect 127711 274961 142857 274989
rect 142885 274961 142919 274989
rect 142947 274961 142981 274989
rect 143009 274961 143043 274989
rect 143071 274961 158217 274989
rect 158245 274961 158279 274989
rect 158307 274961 158341 274989
rect 158369 274961 158403 274989
rect 158431 274961 173577 274989
rect 173605 274961 173639 274989
rect 173667 274961 173701 274989
rect 173729 274961 173763 274989
rect 173791 274961 188937 274989
rect 188965 274961 188999 274989
rect 189027 274961 189061 274989
rect 189089 274961 189123 274989
rect 189151 274961 204297 274989
rect 204325 274961 204359 274989
rect 204387 274961 204421 274989
rect 204449 274961 204483 274989
rect 204511 274961 219657 274989
rect 219685 274961 219719 274989
rect 219747 274961 219781 274989
rect 219809 274961 219843 274989
rect 219871 274961 235017 274989
rect 235045 274961 235079 274989
rect 235107 274961 235141 274989
rect 235169 274961 235203 274989
rect 235231 274961 250377 274989
rect 250405 274961 250439 274989
rect 250467 274961 250501 274989
rect 250529 274961 250563 274989
rect 250591 274961 265737 274989
rect 265765 274961 265799 274989
rect 265827 274961 265861 274989
rect 265889 274961 265923 274989
rect 265951 274961 281097 274989
rect 281125 274961 281159 274989
rect 281187 274961 281221 274989
rect 281249 274961 281283 274989
rect 281311 274961 296457 274989
rect 296485 274961 296519 274989
rect 296547 274961 296581 274989
rect 296609 274961 296643 274989
rect 296671 274961 298728 274989
rect 298756 274961 298790 274989
rect 298818 274961 298852 274989
rect 298880 274961 298914 274989
rect 298942 274961 298990 274989
rect -958 274913 298990 274961
rect -958 272175 298990 272223
rect -958 272147 -430 272175
rect -402 272147 -368 272175
rect -340 272147 -306 272175
rect -278 272147 -244 272175
rect -216 272147 2757 272175
rect 2785 272147 2819 272175
rect 2847 272147 2881 272175
rect 2909 272147 2943 272175
rect 2971 272147 18117 272175
rect 18145 272147 18179 272175
rect 18207 272147 18241 272175
rect 18269 272147 18303 272175
rect 18331 272147 33477 272175
rect 33505 272147 33539 272175
rect 33567 272147 33601 272175
rect 33629 272147 33663 272175
rect 33691 272147 48837 272175
rect 48865 272147 48899 272175
rect 48927 272147 48961 272175
rect 48989 272147 49023 272175
rect 49051 272147 64197 272175
rect 64225 272147 64259 272175
rect 64287 272147 64321 272175
rect 64349 272147 64383 272175
rect 64411 272147 79557 272175
rect 79585 272147 79619 272175
rect 79647 272147 79681 272175
rect 79709 272147 79743 272175
rect 79771 272147 94917 272175
rect 94945 272147 94979 272175
rect 95007 272147 95041 272175
rect 95069 272147 95103 272175
rect 95131 272147 110277 272175
rect 110305 272147 110339 272175
rect 110367 272147 110401 272175
rect 110429 272147 110463 272175
rect 110491 272147 125637 272175
rect 125665 272147 125699 272175
rect 125727 272147 125761 272175
rect 125789 272147 125823 272175
rect 125851 272147 140997 272175
rect 141025 272147 141059 272175
rect 141087 272147 141121 272175
rect 141149 272147 141183 272175
rect 141211 272147 156357 272175
rect 156385 272147 156419 272175
rect 156447 272147 156481 272175
rect 156509 272147 156543 272175
rect 156571 272147 171717 272175
rect 171745 272147 171779 272175
rect 171807 272147 171841 272175
rect 171869 272147 171903 272175
rect 171931 272147 187077 272175
rect 187105 272147 187139 272175
rect 187167 272147 187201 272175
rect 187229 272147 187263 272175
rect 187291 272147 202437 272175
rect 202465 272147 202499 272175
rect 202527 272147 202561 272175
rect 202589 272147 202623 272175
rect 202651 272147 217797 272175
rect 217825 272147 217859 272175
rect 217887 272147 217921 272175
rect 217949 272147 217983 272175
rect 218011 272147 233157 272175
rect 233185 272147 233219 272175
rect 233247 272147 233281 272175
rect 233309 272147 233343 272175
rect 233371 272147 248517 272175
rect 248545 272147 248579 272175
rect 248607 272147 248641 272175
rect 248669 272147 248703 272175
rect 248731 272147 263877 272175
rect 263905 272147 263939 272175
rect 263967 272147 264001 272175
rect 264029 272147 264063 272175
rect 264091 272147 279237 272175
rect 279265 272147 279299 272175
rect 279327 272147 279361 272175
rect 279389 272147 279423 272175
rect 279451 272147 294597 272175
rect 294625 272147 294659 272175
rect 294687 272147 294721 272175
rect 294749 272147 294783 272175
rect 294811 272147 298248 272175
rect 298276 272147 298310 272175
rect 298338 272147 298372 272175
rect 298400 272147 298434 272175
rect 298462 272147 298990 272175
rect -958 272113 298990 272147
rect -958 272085 -430 272113
rect -402 272085 -368 272113
rect -340 272085 -306 272113
rect -278 272085 -244 272113
rect -216 272085 2757 272113
rect 2785 272085 2819 272113
rect 2847 272085 2881 272113
rect 2909 272085 2943 272113
rect 2971 272085 18117 272113
rect 18145 272085 18179 272113
rect 18207 272085 18241 272113
rect 18269 272085 18303 272113
rect 18331 272085 33477 272113
rect 33505 272085 33539 272113
rect 33567 272085 33601 272113
rect 33629 272085 33663 272113
rect 33691 272085 48837 272113
rect 48865 272085 48899 272113
rect 48927 272085 48961 272113
rect 48989 272085 49023 272113
rect 49051 272085 64197 272113
rect 64225 272085 64259 272113
rect 64287 272085 64321 272113
rect 64349 272085 64383 272113
rect 64411 272085 79557 272113
rect 79585 272085 79619 272113
rect 79647 272085 79681 272113
rect 79709 272085 79743 272113
rect 79771 272085 94917 272113
rect 94945 272085 94979 272113
rect 95007 272085 95041 272113
rect 95069 272085 95103 272113
rect 95131 272085 110277 272113
rect 110305 272085 110339 272113
rect 110367 272085 110401 272113
rect 110429 272085 110463 272113
rect 110491 272085 125637 272113
rect 125665 272085 125699 272113
rect 125727 272085 125761 272113
rect 125789 272085 125823 272113
rect 125851 272085 140997 272113
rect 141025 272085 141059 272113
rect 141087 272085 141121 272113
rect 141149 272085 141183 272113
rect 141211 272085 156357 272113
rect 156385 272085 156419 272113
rect 156447 272085 156481 272113
rect 156509 272085 156543 272113
rect 156571 272085 171717 272113
rect 171745 272085 171779 272113
rect 171807 272085 171841 272113
rect 171869 272085 171903 272113
rect 171931 272085 187077 272113
rect 187105 272085 187139 272113
rect 187167 272085 187201 272113
rect 187229 272085 187263 272113
rect 187291 272085 202437 272113
rect 202465 272085 202499 272113
rect 202527 272085 202561 272113
rect 202589 272085 202623 272113
rect 202651 272085 217797 272113
rect 217825 272085 217859 272113
rect 217887 272085 217921 272113
rect 217949 272085 217983 272113
rect 218011 272085 233157 272113
rect 233185 272085 233219 272113
rect 233247 272085 233281 272113
rect 233309 272085 233343 272113
rect 233371 272085 248517 272113
rect 248545 272085 248579 272113
rect 248607 272085 248641 272113
rect 248669 272085 248703 272113
rect 248731 272085 263877 272113
rect 263905 272085 263939 272113
rect 263967 272085 264001 272113
rect 264029 272085 264063 272113
rect 264091 272085 279237 272113
rect 279265 272085 279299 272113
rect 279327 272085 279361 272113
rect 279389 272085 279423 272113
rect 279451 272085 294597 272113
rect 294625 272085 294659 272113
rect 294687 272085 294721 272113
rect 294749 272085 294783 272113
rect 294811 272085 298248 272113
rect 298276 272085 298310 272113
rect 298338 272085 298372 272113
rect 298400 272085 298434 272113
rect 298462 272085 298990 272113
rect -958 272051 298990 272085
rect -958 272023 -430 272051
rect -402 272023 -368 272051
rect -340 272023 -306 272051
rect -278 272023 -244 272051
rect -216 272023 2757 272051
rect 2785 272023 2819 272051
rect 2847 272023 2881 272051
rect 2909 272023 2943 272051
rect 2971 272023 18117 272051
rect 18145 272023 18179 272051
rect 18207 272023 18241 272051
rect 18269 272023 18303 272051
rect 18331 272023 33477 272051
rect 33505 272023 33539 272051
rect 33567 272023 33601 272051
rect 33629 272023 33663 272051
rect 33691 272023 48837 272051
rect 48865 272023 48899 272051
rect 48927 272023 48961 272051
rect 48989 272023 49023 272051
rect 49051 272023 64197 272051
rect 64225 272023 64259 272051
rect 64287 272023 64321 272051
rect 64349 272023 64383 272051
rect 64411 272023 79557 272051
rect 79585 272023 79619 272051
rect 79647 272023 79681 272051
rect 79709 272023 79743 272051
rect 79771 272023 94917 272051
rect 94945 272023 94979 272051
rect 95007 272023 95041 272051
rect 95069 272023 95103 272051
rect 95131 272023 110277 272051
rect 110305 272023 110339 272051
rect 110367 272023 110401 272051
rect 110429 272023 110463 272051
rect 110491 272023 125637 272051
rect 125665 272023 125699 272051
rect 125727 272023 125761 272051
rect 125789 272023 125823 272051
rect 125851 272023 140997 272051
rect 141025 272023 141059 272051
rect 141087 272023 141121 272051
rect 141149 272023 141183 272051
rect 141211 272023 156357 272051
rect 156385 272023 156419 272051
rect 156447 272023 156481 272051
rect 156509 272023 156543 272051
rect 156571 272023 171717 272051
rect 171745 272023 171779 272051
rect 171807 272023 171841 272051
rect 171869 272023 171903 272051
rect 171931 272023 187077 272051
rect 187105 272023 187139 272051
rect 187167 272023 187201 272051
rect 187229 272023 187263 272051
rect 187291 272023 202437 272051
rect 202465 272023 202499 272051
rect 202527 272023 202561 272051
rect 202589 272023 202623 272051
rect 202651 272023 217797 272051
rect 217825 272023 217859 272051
rect 217887 272023 217921 272051
rect 217949 272023 217983 272051
rect 218011 272023 233157 272051
rect 233185 272023 233219 272051
rect 233247 272023 233281 272051
rect 233309 272023 233343 272051
rect 233371 272023 248517 272051
rect 248545 272023 248579 272051
rect 248607 272023 248641 272051
rect 248669 272023 248703 272051
rect 248731 272023 263877 272051
rect 263905 272023 263939 272051
rect 263967 272023 264001 272051
rect 264029 272023 264063 272051
rect 264091 272023 279237 272051
rect 279265 272023 279299 272051
rect 279327 272023 279361 272051
rect 279389 272023 279423 272051
rect 279451 272023 294597 272051
rect 294625 272023 294659 272051
rect 294687 272023 294721 272051
rect 294749 272023 294783 272051
rect 294811 272023 298248 272051
rect 298276 272023 298310 272051
rect 298338 272023 298372 272051
rect 298400 272023 298434 272051
rect 298462 272023 298990 272051
rect -958 271989 298990 272023
rect -958 271961 -430 271989
rect -402 271961 -368 271989
rect -340 271961 -306 271989
rect -278 271961 -244 271989
rect -216 271961 2757 271989
rect 2785 271961 2819 271989
rect 2847 271961 2881 271989
rect 2909 271961 2943 271989
rect 2971 271961 18117 271989
rect 18145 271961 18179 271989
rect 18207 271961 18241 271989
rect 18269 271961 18303 271989
rect 18331 271961 33477 271989
rect 33505 271961 33539 271989
rect 33567 271961 33601 271989
rect 33629 271961 33663 271989
rect 33691 271961 48837 271989
rect 48865 271961 48899 271989
rect 48927 271961 48961 271989
rect 48989 271961 49023 271989
rect 49051 271961 64197 271989
rect 64225 271961 64259 271989
rect 64287 271961 64321 271989
rect 64349 271961 64383 271989
rect 64411 271961 79557 271989
rect 79585 271961 79619 271989
rect 79647 271961 79681 271989
rect 79709 271961 79743 271989
rect 79771 271961 94917 271989
rect 94945 271961 94979 271989
rect 95007 271961 95041 271989
rect 95069 271961 95103 271989
rect 95131 271961 110277 271989
rect 110305 271961 110339 271989
rect 110367 271961 110401 271989
rect 110429 271961 110463 271989
rect 110491 271961 125637 271989
rect 125665 271961 125699 271989
rect 125727 271961 125761 271989
rect 125789 271961 125823 271989
rect 125851 271961 140997 271989
rect 141025 271961 141059 271989
rect 141087 271961 141121 271989
rect 141149 271961 141183 271989
rect 141211 271961 156357 271989
rect 156385 271961 156419 271989
rect 156447 271961 156481 271989
rect 156509 271961 156543 271989
rect 156571 271961 171717 271989
rect 171745 271961 171779 271989
rect 171807 271961 171841 271989
rect 171869 271961 171903 271989
rect 171931 271961 187077 271989
rect 187105 271961 187139 271989
rect 187167 271961 187201 271989
rect 187229 271961 187263 271989
rect 187291 271961 202437 271989
rect 202465 271961 202499 271989
rect 202527 271961 202561 271989
rect 202589 271961 202623 271989
rect 202651 271961 217797 271989
rect 217825 271961 217859 271989
rect 217887 271961 217921 271989
rect 217949 271961 217983 271989
rect 218011 271961 233157 271989
rect 233185 271961 233219 271989
rect 233247 271961 233281 271989
rect 233309 271961 233343 271989
rect 233371 271961 248517 271989
rect 248545 271961 248579 271989
rect 248607 271961 248641 271989
rect 248669 271961 248703 271989
rect 248731 271961 263877 271989
rect 263905 271961 263939 271989
rect 263967 271961 264001 271989
rect 264029 271961 264063 271989
rect 264091 271961 279237 271989
rect 279265 271961 279299 271989
rect 279327 271961 279361 271989
rect 279389 271961 279423 271989
rect 279451 271961 294597 271989
rect 294625 271961 294659 271989
rect 294687 271961 294721 271989
rect 294749 271961 294783 271989
rect 294811 271961 298248 271989
rect 298276 271961 298310 271989
rect 298338 271961 298372 271989
rect 298400 271961 298434 271989
rect 298462 271961 298990 271989
rect -958 271913 298990 271961
rect -958 266175 298990 266223
rect -958 266147 -910 266175
rect -882 266147 -848 266175
rect -820 266147 -786 266175
rect -758 266147 -724 266175
rect -696 266147 4617 266175
rect 4645 266147 4679 266175
rect 4707 266147 4741 266175
rect 4769 266147 4803 266175
rect 4831 266147 29939 266175
rect 29967 266147 30001 266175
rect 30029 266147 45299 266175
rect 45327 266147 45361 266175
rect 45389 266147 60659 266175
rect 60687 266147 60721 266175
rect 60749 266147 76019 266175
rect 76047 266147 76081 266175
rect 76109 266147 96777 266175
rect 96805 266147 96839 266175
rect 96867 266147 96901 266175
rect 96929 266147 96963 266175
rect 96991 266147 109939 266175
rect 109967 266147 110001 266175
rect 110029 266147 125299 266175
rect 125327 266147 125361 266175
rect 125389 266147 140659 266175
rect 140687 266147 140721 266175
rect 140749 266147 156019 266175
rect 156047 266147 156081 266175
rect 156109 266147 173577 266175
rect 173605 266147 173639 266175
rect 173667 266147 173701 266175
rect 173729 266147 173763 266175
rect 173791 266147 188937 266175
rect 188965 266147 188999 266175
rect 189027 266147 189061 266175
rect 189089 266147 189123 266175
rect 189151 266147 204297 266175
rect 204325 266147 204359 266175
rect 204387 266147 204421 266175
rect 204449 266147 204483 266175
rect 204511 266147 219657 266175
rect 219685 266147 219719 266175
rect 219747 266147 219781 266175
rect 219809 266147 219843 266175
rect 219871 266147 235017 266175
rect 235045 266147 235079 266175
rect 235107 266147 235141 266175
rect 235169 266147 235203 266175
rect 235231 266147 250377 266175
rect 250405 266147 250439 266175
rect 250467 266147 250501 266175
rect 250529 266147 250563 266175
rect 250591 266147 265737 266175
rect 265765 266147 265799 266175
rect 265827 266147 265861 266175
rect 265889 266147 265923 266175
rect 265951 266147 281097 266175
rect 281125 266147 281159 266175
rect 281187 266147 281221 266175
rect 281249 266147 281283 266175
rect 281311 266147 296457 266175
rect 296485 266147 296519 266175
rect 296547 266147 296581 266175
rect 296609 266147 296643 266175
rect 296671 266147 298728 266175
rect 298756 266147 298790 266175
rect 298818 266147 298852 266175
rect 298880 266147 298914 266175
rect 298942 266147 298990 266175
rect -958 266113 298990 266147
rect -958 266085 -910 266113
rect -882 266085 -848 266113
rect -820 266085 -786 266113
rect -758 266085 -724 266113
rect -696 266085 4617 266113
rect 4645 266085 4679 266113
rect 4707 266085 4741 266113
rect 4769 266085 4803 266113
rect 4831 266085 29939 266113
rect 29967 266085 30001 266113
rect 30029 266085 45299 266113
rect 45327 266085 45361 266113
rect 45389 266085 60659 266113
rect 60687 266085 60721 266113
rect 60749 266085 76019 266113
rect 76047 266085 76081 266113
rect 76109 266085 96777 266113
rect 96805 266085 96839 266113
rect 96867 266085 96901 266113
rect 96929 266085 96963 266113
rect 96991 266085 109939 266113
rect 109967 266085 110001 266113
rect 110029 266085 125299 266113
rect 125327 266085 125361 266113
rect 125389 266085 140659 266113
rect 140687 266085 140721 266113
rect 140749 266085 156019 266113
rect 156047 266085 156081 266113
rect 156109 266085 173577 266113
rect 173605 266085 173639 266113
rect 173667 266085 173701 266113
rect 173729 266085 173763 266113
rect 173791 266085 188937 266113
rect 188965 266085 188999 266113
rect 189027 266085 189061 266113
rect 189089 266085 189123 266113
rect 189151 266085 204297 266113
rect 204325 266085 204359 266113
rect 204387 266085 204421 266113
rect 204449 266085 204483 266113
rect 204511 266085 219657 266113
rect 219685 266085 219719 266113
rect 219747 266085 219781 266113
rect 219809 266085 219843 266113
rect 219871 266085 235017 266113
rect 235045 266085 235079 266113
rect 235107 266085 235141 266113
rect 235169 266085 235203 266113
rect 235231 266085 250377 266113
rect 250405 266085 250439 266113
rect 250467 266085 250501 266113
rect 250529 266085 250563 266113
rect 250591 266085 265737 266113
rect 265765 266085 265799 266113
rect 265827 266085 265861 266113
rect 265889 266085 265923 266113
rect 265951 266085 281097 266113
rect 281125 266085 281159 266113
rect 281187 266085 281221 266113
rect 281249 266085 281283 266113
rect 281311 266085 296457 266113
rect 296485 266085 296519 266113
rect 296547 266085 296581 266113
rect 296609 266085 296643 266113
rect 296671 266085 298728 266113
rect 298756 266085 298790 266113
rect 298818 266085 298852 266113
rect 298880 266085 298914 266113
rect 298942 266085 298990 266113
rect -958 266051 298990 266085
rect -958 266023 -910 266051
rect -882 266023 -848 266051
rect -820 266023 -786 266051
rect -758 266023 -724 266051
rect -696 266023 4617 266051
rect 4645 266023 4679 266051
rect 4707 266023 4741 266051
rect 4769 266023 4803 266051
rect 4831 266023 29939 266051
rect 29967 266023 30001 266051
rect 30029 266023 45299 266051
rect 45327 266023 45361 266051
rect 45389 266023 60659 266051
rect 60687 266023 60721 266051
rect 60749 266023 76019 266051
rect 76047 266023 76081 266051
rect 76109 266023 96777 266051
rect 96805 266023 96839 266051
rect 96867 266023 96901 266051
rect 96929 266023 96963 266051
rect 96991 266023 109939 266051
rect 109967 266023 110001 266051
rect 110029 266023 125299 266051
rect 125327 266023 125361 266051
rect 125389 266023 140659 266051
rect 140687 266023 140721 266051
rect 140749 266023 156019 266051
rect 156047 266023 156081 266051
rect 156109 266023 173577 266051
rect 173605 266023 173639 266051
rect 173667 266023 173701 266051
rect 173729 266023 173763 266051
rect 173791 266023 188937 266051
rect 188965 266023 188999 266051
rect 189027 266023 189061 266051
rect 189089 266023 189123 266051
rect 189151 266023 204297 266051
rect 204325 266023 204359 266051
rect 204387 266023 204421 266051
rect 204449 266023 204483 266051
rect 204511 266023 219657 266051
rect 219685 266023 219719 266051
rect 219747 266023 219781 266051
rect 219809 266023 219843 266051
rect 219871 266023 235017 266051
rect 235045 266023 235079 266051
rect 235107 266023 235141 266051
rect 235169 266023 235203 266051
rect 235231 266023 250377 266051
rect 250405 266023 250439 266051
rect 250467 266023 250501 266051
rect 250529 266023 250563 266051
rect 250591 266023 265737 266051
rect 265765 266023 265799 266051
rect 265827 266023 265861 266051
rect 265889 266023 265923 266051
rect 265951 266023 281097 266051
rect 281125 266023 281159 266051
rect 281187 266023 281221 266051
rect 281249 266023 281283 266051
rect 281311 266023 296457 266051
rect 296485 266023 296519 266051
rect 296547 266023 296581 266051
rect 296609 266023 296643 266051
rect 296671 266023 298728 266051
rect 298756 266023 298790 266051
rect 298818 266023 298852 266051
rect 298880 266023 298914 266051
rect 298942 266023 298990 266051
rect -958 265989 298990 266023
rect -958 265961 -910 265989
rect -882 265961 -848 265989
rect -820 265961 -786 265989
rect -758 265961 -724 265989
rect -696 265961 4617 265989
rect 4645 265961 4679 265989
rect 4707 265961 4741 265989
rect 4769 265961 4803 265989
rect 4831 265961 29939 265989
rect 29967 265961 30001 265989
rect 30029 265961 45299 265989
rect 45327 265961 45361 265989
rect 45389 265961 60659 265989
rect 60687 265961 60721 265989
rect 60749 265961 76019 265989
rect 76047 265961 76081 265989
rect 76109 265961 96777 265989
rect 96805 265961 96839 265989
rect 96867 265961 96901 265989
rect 96929 265961 96963 265989
rect 96991 265961 109939 265989
rect 109967 265961 110001 265989
rect 110029 265961 125299 265989
rect 125327 265961 125361 265989
rect 125389 265961 140659 265989
rect 140687 265961 140721 265989
rect 140749 265961 156019 265989
rect 156047 265961 156081 265989
rect 156109 265961 173577 265989
rect 173605 265961 173639 265989
rect 173667 265961 173701 265989
rect 173729 265961 173763 265989
rect 173791 265961 188937 265989
rect 188965 265961 188999 265989
rect 189027 265961 189061 265989
rect 189089 265961 189123 265989
rect 189151 265961 204297 265989
rect 204325 265961 204359 265989
rect 204387 265961 204421 265989
rect 204449 265961 204483 265989
rect 204511 265961 219657 265989
rect 219685 265961 219719 265989
rect 219747 265961 219781 265989
rect 219809 265961 219843 265989
rect 219871 265961 235017 265989
rect 235045 265961 235079 265989
rect 235107 265961 235141 265989
rect 235169 265961 235203 265989
rect 235231 265961 250377 265989
rect 250405 265961 250439 265989
rect 250467 265961 250501 265989
rect 250529 265961 250563 265989
rect 250591 265961 265737 265989
rect 265765 265961 265799 265989
rect 265827 265961 265861 265989
rect 265889 265961 265923 265989
rect 265951 265961 281097 265989
rect 281125 265961 281159 265989
rect 281187 265961 281221 265989
rect 281249 265961 281283 265989
rect 281311 265961 296457 265989
rect 296485 265961 296519 265989
rect 296547 265961 296581 265989
rect 296609 265961 296643 265989
rect 296671 265961 298728 265989
rect 298756 265961 298790 265989
rect 298818 265961 298852 265989
rect 298880 265961 298914 265989
rect 298942 265961 298990 265989
rect -958 265913 298990 265961
rect -958 263175 298990 263223
rect -958 263147 -430 263175
rect -402 263147 -368 263175
rect -340 263147 -306 263175
rect -278 263147 -244 263175
rect -216 263147 2757 263175
rect 2785 263147 2819 263175
rect 2847 263147 2881 263175
rect 2909 263147 2943 263175
rect 2971 263147 18117 263175
rect 18145 263147 18179 263175
rect 18207 263147 18241 263175
rect 18269 263147 18303 263175
rect 18331 263147 22259 263175
rect 22287 263147 22321 263175
rect 22349 263147 37619 263175
rect 37647 263147 37681 263175
rect 37709 263147 52979 263175
rect 53007 263147 53041 263175
rect 53069 263147 68339 263175
rect 68367 263147 68401 263175
rect 68429 263147 83699 263175
rect 83727 263147 83761 263175
rect 83789 263147 94917 263175
rect 94945 263147 94979 263175
rect 95007 263147 95041 263175
rect 95069 263147 95103 263175
rect 95131 263147 102259 263175
rect 102287 263147 102321 263175
rect 102349 263147 117619 263175
rect 117647 263147 117681 263175
rect 117709 263147 132979 263175
rect 133007 263147 133041 263175
rect 133069 263147 148339 263175
rect 148367 263147 148401 263175
rect 148429 263147 163699 263175
rect 163727 263147 163761 263175
rect 163789 263147 171717 263175
rect 171745 263147 171779 263175
rect 171807 263147 171841 263175
rect 171869 263147 171903 263175
rect 171931 263147 187077 263175
rect 187105 263147 187139 263175
rect 187167 263147 187201 263175
rect 187229 263147 187263 263175
rect 187291 263147 202437 263175
rect 202465 263147 202499 263175
rect 202527 263147 202561 263175
rect 202589 263147 202623 263175
rect 202651 263147 217797 263175
rect 217825 263147 217859 263175
rect 217887 263147 217921 263175
rect 217949 263147 217983 263175
rect 218011 263147 233157 263175
rect 233185 263147 233219 263175
rect 233247 263147 233281 263175
rect 233309 263147 233343 263175
rect 233371 263147 248517 263175
rect 248545 263147 248579 263175
rect 248607 263147 248641 263175
rect 248669 263147 248703 263175
rect 248731 263147 263877 263175
rect 263905 263147 263939 263175
rect 263967 263147 264001 263175
rect 264029 263147 264063 263175
rect 264091 263147 279237 263175
rect 279265 263147 279299 263175
rect 279327 263147 279361 263175
rect 279389 263147 279423 263175
rect 279451 263147 294597 263175
rect 294625 263147 294659 263175
rect 294687 263147 294721 263175
rect 294749 263147 294783 263175
rect 294811 263147 298248 263175
rect 298276 263147 298310 263175
rect 298338 263147 298372 263175
rect 298400 263147 298434 263175
rect 298462 263147 298990 263175
rect -958 263113 298990 263147
rect -958 263085 -430 263113
rect -402 263085 -368 263113
rect -340 263085 -306 263113
rect -278 263085 -244 263113
rect -216 263085 2757 263113
rect 2785 263085 2819 263113
rect 2847 263085 2881 263113
rect 2909 263085 2943 263113
rect 2971 263085 18117 263113
rect 18145 263085 18179 263113
rect 18207 263085 18241 263113
rect 18269 263085 18303 263113
rect 18331 263085 22259 263113
rect 22287 263085 22321 263113
rect 22349 263085 37619 263113
rect 37647 263085 37681 263113
rect 37709 263085 52979 263113
rect 53007 263085 53041 263113
rect 53069 263085 68339 263113
rect 68367 263085 68401 263113
rect 68429 263085 83699 263113
rect 83727 263085 83761 263113
rect 83789 263085 94917 263113
rect 94945 263085 94979 263113
rect 95007 263085 95041 263113
rect 95069 263085 95103 263113
rect 95131 263085 102259 263113
rect 102287 263085 102321 263113
rect 102349 263085 117619 263113
rect 117647 263085 117681 263113
rect 117709 263085 132979 263113
rect 133007 263085 133041 263113
rect 133069 263085 148339 263113
rect 148367 263085 148401 263113
rect 148429 263085 163699 263113
rect 163727 263085 163761 263113
rect 163789 263085 171717 263113
rect 171745 263085 171779 263113
rect 171807 263085 171841 263113
rect 171869 263085 171903 263113
rect 171931 263085 187077 263113
rect 187105 263085 187139 263113
rect 187167 263085 187201 263113
rect 187229 263085 187263 263113
rect 187291 263085 202437 263113
rect 202465 263085 202499 263113
rect 202527 263085 202561 263113
rect 202589 263085 202623 263113
rect 202651 263085 217797 263113
rect 217825 263085 217859 263113
rect 217887 263085 217921 263113
rect 217949 263085 217983 263113
rect 218011 263085 233157 263113
rect 233185 263085 233219 263113
rect 233247 263085 233281 263113
rect 233309 263085 233343 263113
rect 233371 263085 248517 263113
rect 248545 263085 248579 263113
rect 248607 263085 248641 263113
rect 248669 263085 248703 263113
rect 248731 263085 263877 263113
rect 263905 263085 263939 263113
rect 263967 263085 264001 263113
rect 264029 263085 264063 263113
rect 264091 263085 279237 263113
rect 279265 263085 279299 263113
rect 279327 263085 279361 263113
rect 279389 263085 279423 263113
rect 279451 263085 294597 263113
rect 294625 263085 294659 263113
rect 294687 263085 294721 263113
rect 294749 263085 294783 263113
rect 294811 263085 298248 263113
rect 298276 263085 298310 263113
rect 298338 263085 298372 263113
rect 298400 263085 298434 263113
rect 298462 263085 298990 263113
rect -958 263051 298990 263085
rect -958 263023 -430 263051
rect -402 263023 -368 263051
rect -340 263023 -306 263051
rect -278 263023 -244 263051
rect -216 263023 2757 263051
rect 2785 263023 2819 263051
rect 2847 263023 2881 263051
rect 2909 263023 2943 263051
rect 2971 263023 18117 263051
rect 18145 263023 18179 263051
rect 18207 263023 18241 263051
rect 18269 263023 18303 263051
rect 18331 263023 22259 263051
rect 22287 263023 22321 263051
rect 22349 263023 37619 263051
rect 37647 263023 37681 263051
rect 37709 263023 52979 263051
rect 53007 263023 53041 263051
rect 53069 263023 68339 263051
rect 68367 263023 68401 263051
rect 68429 263023 83699 263051
rect 83727 263023 83761 263051
rect 83789 263023 94917 263051
rect 94945 263023 94979 263051
rect 95007 263023 95041 263051
rect 95069 263023 95103 263051
rect 95131 263023 102259 263051
rect 102287 263023 102321 263051
rect 102349 263023 117619 263051
rect 117647 263023 117681 263051
rect 117709 263023 132979 263051
rect 133007 263023 133041 263051
rect 133069 263023 148339 263051
rect 148367 263023 148401 263051
rect 148429 263023 163699 263051
rect 163727 263023 163761 263051
rect 163789 263023 171717 263051
rect 171745 263023 171779 263051
rect 171807 263023 171841 263051
rect 171869 263023 171903 263051
rect 171931 263023 187077 263051
rect 187105 263023 187139 263051
rect 187167 263023 187201 263051
rect 187229 263023 187263 263051
rect 187291 263023 202437 263051
rect 202465 263023 202499 263051
rect 202527 263023 202561 263051
rect 202589 263023 202623 263051
rect 202651 263023 217797 263051
rect 217825 263023 217859 263051
rect 217887 263023 217921 263051
rect 217949 263023 217983 263051
rect 218011 263023 233157 263051
rect 233185 263023 233219 263051
rect 233247 263023 233281 263051
rect 233309 263023 233343 263051
rect 233371 263023 248517 263051
rect 248545 263023 248579 263051
rect 248607 263023 248641 263051
rect 248669 263023 248703 263051
rect 248731 263023 263877 263051
rect 263905 263023 263939 263051
rect 263967 263023 264001 263051
rect 264029 263023 264063 263051
rect 264091 263023 279237 263051
rect 279265 263023 279299 263051
rect 279327 263023 279361 263051
rect 279389 263023 279423 263051
rect 279451 263023 294597 263051
rect 294625 263023 294659 263051
rect 294687 263023 294721 263051
rect 294749 263023 294783 263051
rect 294811 263023 298248 263051
rect 298276 263023 298310 263051
rect 298338 263023 298372 263051
rect 298400 263023 298434 263051
rect 298462 263023 298990 263051
rect -958 262989 298990 263023
rect -958 262961 -430 262989
rect -402 262961 -368 262989
rect -340 262961 -306 262989
rect -278 262961 -244 262989
rect -216 262961 2757 262989
rect 2785 262961 2819 262989
rect 2847 262961 2881 262989
rect 2909 262961 2943 262989
rect 2971 262961 18117 262989
rect 18145 262961 18179 262989
rect 18207 262961 18241 262989
rect 18269 262961 18303 262989
rect 18331 262961 22259 262989
rect 22287 262961 22321 262989
rect 22349 262961 37619 262989
rect 37647 262961 37681 262989
rect 37709 262961 52979 262989
rect 53007 262961 53041 262989
rect 53069 262961 68339 262989
rect 68367 262961 68401 262989
rect 68429 262961 83699 262989
rect 83727 262961 83761 262989
rect 83789 262961 94917 262989
rect 94945 262961 94979 262989
rect 95007 262961 95041 262989
rect 95069 262961 95103 262989
rect 95131 262961 102259 262989
rect 102287 262961 102321 262989
rect 102349 262961 117619 262989
rect 117647 262961 117681 262989
rect 117709 262961 132979 262989
rect 133007 262961 133041 262989
rect 133069 262961 148339 262989
rect 148367 262961 148401 262989
rect 148429 262961 163699 262989
rect 163727 262961 163761 262989
rect 163789 262961 171717 262989
rect 171745 262961 171779 262989
rect 171807 262961 171841 262989
rect 171869 262961 171903 262989
rect 171931 262961 187077 262989
rect 187105 262961 187139 262989
rect 187167 262961 187201 262989
rect 187229 262961 187263 262989
rect 187291 262961 202437 262989
rect 202465 262961 202499 262989
rect 202527 262961 202561 262989
rect 202589 262961 202623 262989
rect 202651 262961 217797 262989
rect 217825 262961 217859 262989
rect 217887 262961 217921 262989
rect 217949 262961 217983 262989
rect 218011 262961 233157 262989
rect 233185 262961 233219 262989
rect 233247 262961 233281 262989
rect 233309 262961 233343 262989
rect 233371 262961 248517 262989
rect 248545 262961 248579 262989
rect 248607 262961 248641 262989
rect 248669 262961 248703 262989
rect 248731 262961 263877 262989
rect 263905 262961 263939 262989
rect 263967 262961 264001 262989
rect 264029 262961 264063 262989
rect 264091 262961 279237 262989
rect 279265 262961 279299 262989
rect 279327 262961 279361 262989
rect 279389 262961 279423 262989
rect 279451 262961 294597 262989
rect 294625 262961 294659 262989
rect 294687 262961 294721 262989
rect 294749 262961 294783 262989
rect 294811 262961 298248 262989
rect 298276 262961 298310 262989
rect 298338 262961 298372 262989
rect 298400 262961 298434 262989
rect 298462 262961 298990 262989
rect -958 262913 298990 262961
rect -958 257175 298990 257223
rect -958 257147 -910 257175
rect -882 257147 -848 257175
rect -820 257147 -786 257175
rect -758 257147 -724 257175
rect -696 257147 4617 257175
rect 4645 257147 4679 257175
rect 4707 257147 4741 257175
rect 4769 257147 4803 257175
rect 4831 257147 29939 257175
rect 29967 257147 30001 257175
rect 30029 257147 45299 257175
rect 45327 257147 45361 257175
rect 45389 257147 60659 257175
rect 60687 257147 60721 257175
rect 60749 257147 76019 257175
rect 76047 257147 76081 257175
rect 76109 257147 96777 257175
rect 96805 257147 96839 257175
rect 96867 257147 96901 257175
rect 96929 257147 96963 257175
rect 96991 257147 109939 257175
rect 109967 257147 110001 257175
rect 110029 257147 125299 257175
rect 125327 257147 125361 257175
rect 125389 257147 140659 257175
rect 140687 257147 140721 257175
rect 140749 257147 156019 257175
rect 156047 257147 156081 257175
rect 156109 257147 173577 257175
rect 173605 257147 173639 257175
rect 173667 257147 173701 257175
rect 173729 257147 173763 257175
rect 173791 257147 188937 257175
rect 188965 257147 188999 257175
rect 189027 257147 189061 257175
rect 189089 257147 189123 257175
rect 189151 257147 204297 257175
rect 204325 257147 204359 257175
rect 204387 257147 204421 257175
rect 204449 257147 204483 257175
rect 204511 257147 219657 257175
rect 219685 257147 219719 257175
rect 219747 257147 219781 257175
rect 219809 257147 219843 257175
rect 219871 257147 235017 257175
rect 235045 257147 235079 257175
rect 235107 257147 235141 257175
rect 235169 257147 235203 257175
rect 235231 257147 250377 257175
rect 250405 257147 250439 257175
rect 250467 257147 250501 257175
rect 250529 257147 250563 257175
rect 250591 257147 265737 257175
rect 265765 257147 265799 257175
rect 265827 257147 265861 257175
rect 265889 257147 265923 257175
rect 265951 257147 281097 257175
rect 281125 257147 281159 257175
rect 281187 257147 281221 257175
rect 281249 257147 281283 257175
rect 281311 257147 296457 257175
rect 296485 257147 296519 257175
rect 296547 257147 296581 257175
rect 296609 257147 296643 257175
rect 296671 257147 298728 257175
rect 298756 257147 298790 257175
rect 298818 257147 298852 257175
rect 298880 257147 298914 257175
rect 298942 257147 298990 257175
rect -958 257113 298990 257147
rect -958 257085 -910 257113
rect -882 257085 -848 257113
rect -820 257085 -786 257113
rect -758 257085 -724 257113
rect -696 257085 4617 257113
rect 4645 257085 4679 257113
rect 4707 257085 4741 257113
rect 4769 257085 4803 257113
rect 4831 257085 29939 257113
rect 29967 257085 30001 257113
rect 30029 257085 45299 257113
rect 45327 257085 45361 257113
rect 45389 257085 60659 257113
rect 60687 257085 60721 257113
rect 60749 257085 76019 257113
rect 76047 257085 76081 257113
rect 76109 257085 96777 257113
rect 96805 257085 96839 257113
rect 96867 257085 96901 257113
rect 96929 257085 96963 257113
rect 96991 257085 109939 257113
rect 109967 257085 110001 257113
rect 110029 257085 125299 257113
rect 125327 257085 125361 257113
rect 125389 257085 140659 257113
rect 140687 257085 140721 257113
rect 140749 257085 156019 257113
rect 156047 257085 156081 257113
rect 156109 257085 173577 257113
rect 173605 257085 173639 257113
rect 173667 257085 173701 257113
rect 173729 257085 173763 257113
rect 173791 257085 188937 257113
rect 188965 257085 188999 257113
rect 189027 257085 189061 257113
rect 189089 257085 189123 257113
rect 189151 257085 204297 257113
rect 204325 257085 204359 257113
rect 204387 257085 204421 257113
rect 204449 257085 204483 257113
rect 204511 257085 219657 257113
rect 219685 257085 219719 257113
rect 219747 257085 219781 257113
rect 219809 257085 219843 257113
rect 219871 257085 235017 257113
rect 235045 257085 235079 257113
rect 235107 257085 235141 257113
rect 235169 257085 235203 257113
rect 235231 257085 250377 257113
rect 250405 257085 250439 257113
rect 250467 257085 250501 257113
rect 250529 257085 250563 257113
rect 250591 257085 265737 257113
rect 265765 257085 265799 257113
rect 265827 257085 265861 257113
rect 265889 257085 265923 257113
rect 265951 257085 281097 257113
rect 281125 257085 281159 257113
rect 281187 257085 281221 257113
rect 281249 257085 281283 257113
rect 281311 257085 296457 257113
rect 296485 257085 296519 257113
rect 296547 257085 296581 257113
rect 296609 257085 296643 257113
rect 296671 257085 298728 257113
rect 298756 257085 298790 257113
rect 298818 257085 298852 257113
rect 298880 257085 298914 257113
rect 298942 257085 298990 257113
rect -958 257051 298990 257085
rect -958 257023 -910 257051
rect -882 257023 -848 257051
rect -820 257023 -786 257051
rect -758 257023 -724 257051
rect -696 257023 4617 257051
rect 4645 257023 4679 257051
rect 4707 257023 4741 257051
rect 4769 257023 4803 257051
rect 4831 257023 29939 257051
rect 29967 257023 30001 257051
rect 30029 257023 45299 257051
rect 45327 257023 45361 257051
rect 45389 257023 60659 257051
rect 60687 257023 60721 257051
rect 60749 257023 76019 257051
rect 76047 257023 76081 257051
rect 76109 257023 96777 257051
rect 96805 257023 96839 257051
rect 96867 257023 96901 257051
rect 96929 257023 96963 257051
rect 96991 257023 109939 257051
rect 109967 257023 110001 257051
rect 110029 257023 125299 257051
rect 125327 257023 125361 257051
rect 125389 257023 140659 257051
rect 140687 257023 140721 257051
rect 140749 257023 156019 257051
rect 156047 257023 156081 257051
rect 156109 257023 173577 257051
rect 173605 257023 173639 257051
rect 173667 257023 173701 257051
rect 173729 257023 173763 257051
rect 173791 257023 188937 257051
rect 188965 257023 188999 257051
rect 189027 257023 189061 257051
rect 189089 257023 189123 257051
rect 189151 257023 204297 257051
rect 204325 257023 204359 257051
rect 204387 257023 204421 257051
rect 204449 257023 204483 257051
rect 204511 257023 219657 257051
rect 219685 257023 219719 257051
rect 219747 257023 219781 257051
rect 219809 257023 219843 257051
rect 219871 257023 235017 257051
rect 235045 257023 235079 257051
rect 235107 257023 235141 257051
rect 235169 257023 235203 257051
rect 235231 257023 250377 257051
rect 250405 257023 250439 257051
rect 250467 257023 250501 257051
rect 250529 257023 250563 257051
rect 250591 257023 265737 257051
rect 265765 257023 265799 257051
rect 265827 257023 265861 257051
rect 265889 257023 265923 257051
rect 265951 257023 281097 257051
rect 281125 257023 281159 257051
rect 281187 257023 281221 257051
rect 281249 257023 281283 257051
rect 281311 257023 296457 257051
rect 296485 257023 296519 257051
rect 296547 257023 296581 257051
rect 296609 257023 296643 257051
rect 296671 257023 298728 257051
rect 298756 257023 298790 257051
rect 298818 257023 298852 257051
rect 298880 257023 298914 257051
rect 298942 257023 298990 257051
rect -958 256989 298990 257023
rect -958 256961 -910 256989
rect -882 256961 -848 256989
rect -820 256961 -786 256989
rect -758 256961 -724 256989
rect -696 256961 4617 256989
rect 4645 256961 4679 256989
rect 4707 256961 4741 256989
rect 4769 256961 4803 256989
rect 4831 256961 29939 256989
rect 29967 256961 30001 256989
rect 30029 256961 45299 256989
rect 45327 256961 45361 256989
rect 45389 256961 60659 256989
rect 60687 256961 60721 256989
rect 60749 256961 76019 256989
rect 76047 256961 76081 256989
rect 76109 256961 96777 256989
rect 96805 256961 96839 256989
rect 96867 256961 96901 256989
rect 96929 256961 96963 256989
rect 96991 256961 109939 256989
rect 109967 256961 110001 256989
rect 110029 256961 125299 256989
rect 125327 256961 125361 256989
rect 125389 256961 140659 256989
rect 140687 256961 140721 256989
rect 140749 256961 156019 256989
rect 156047 256961 156081 256989
rect 156109 256961 173577 256989
rect 173605 256961 173639 256989
rect 173667 256961 173701 256989
rect 173729 256961 173763 256989
rect 173791 256961 188937 256989
rect 188965 256961 188999 256989
rect 189027 256961 189061 256989
rect 189089 256961 189123 256989
rect 189151 256961 204297 256989
rect 204325 256961 204359 256989
rect 204387 256961 204421 256989
rect 204449 256961 204483 256989
rect 204511 256961 219657 256989
rect 219685 256961 219719 256989
rect 219747 256961 219781 256989
rect 219809 256961 219843 256989
rect 219871 256961 235017 256989
rect 235045 256961 235079 256989
rect 235107 256961 235141 256989
rect 235169 256961 235203 256989
rect 235231 256961 250377 256989
rect 250405 256961 250439 256989
rect 250467 256961 250501 256989
rect 250529 256961 250563 256989
rect 250591 256961 265737 256989
rect 265765 256961 265799 256989
rect 265827 256961 265861 256989
rect 265889 256961 265923 256989
rect 265951 256961 281097 256989
rect 281125 256961 281159 256989
rect 281187 256961 281221 256989
rect 281249 256961 281283 256989
rect 281311 256961 296457 256989
rect 296485 256961 296519 256989
rect 296547 256961 296581 256989
rect 296609 256961 296643 256989
rect 296671 256961 298728 256989
rect 298756 256961 298790 256989
rect 298818 256961 298852 256989
rect 298880 256961 298914 256989
rect 298942 256961 298990 256989
rect -958 256913 298990 256961
rect -958 254175 298990 254223
rect -958 254147 -430 254175
rect -402 254147 -368 254175
rect -340 254147 -306 254175
rect -278 254147 -244 254175
rect -216 254147 2757 254175
rect 2785 254147 2819 254175
rect 2847 254147 2881 254175
rect 2909 254147 2943 254175
rect 2971 254147 18117 254175
rect 18145 254147 18179 254175
rect 18207 254147 18241 254175
rect 18269 254147 18303 254175
rect 18331 254147 22259 254175
rect 22287 254147 22321 254175
rect 22349 254147 37619 254175
rect 37647 254147 37681 254175
rect 37709 254147 52979 254175
rect 53007 254147 53041 254175
rect 53069 254147 68339 254175
rect 68367 254147 68401 254175
rect 68429 254147 83699 254175
rect 83727 254147 83761 254175
rect 83789 254147 94917 254175
rect 94945 254147 94979 254175
rect 95007 254147 95041 254175
rect 95069 254147 95103 254175
rect 95131 254147 102259 254175
rect 102287 254147 102321 254175
rect 102349 254147 117619 254175
rect 117647 254147 117681 254175
rect 117709 254147 132979 254175
rect 133007 254147 133041 254175
rect 133069 254147 148339 254175
rect 148367 254147 148401 254175
rect 148429 254147 163699 254175
rect 163727 254147 163761 254175
rect 163789 254147 171717 254175
rect 171745 254147 171779 254175
rect 171807 254147 171841 254175
rect 171869 254147 171903 254175
rect 171931 254147 187077 254175
rect 187105 254147 187139 254175
rect 187167 254147 187201 254175
rect 187229 254147 187263 254175
rect 187291 254147 202437 254175
rect 202465 254147 202499 254175
rect 202527 254147 202561 254175
rect 202589 254147 202623 254175
rect 202651 254147 217797 254175
rect 217825 254147 217859 254175
rect 217887 254147 217921 254175
rect 217949 254147 217983 254175
rect 218011 254147 233157 254175
rect 233185 254147 233219 254175
rect 233247 254147 233281 254175
rect 233309 254147 233343 254175
rect 233371 254147 248517 254175
rect 248545 254147 248579 254175
rect 248607 254147 248641 254175
rect 248669 254147 248703 254175
rect 248731 254147 263877 254175
rect 263905 254147 263939 254175
rect 263967 254147 264001 254175
rect 264029 254147 264063 254175
rect 264091 254147 279237 254175
rect 279265 254147 279299 254175
rect 279327 254147 279361 254175
rect 279389 254147 279423 254175
rect 279451 254147 294597 254175
rect 294625 254147 294659 254175
rect 294687 254147 294721 254175
rect 294749 254147 294783 254175
rect 294811 254147 298248 254175
rect 298276 254147 298310 254175
rect 298338 254147 298372 254175
rect 298400 254147 298434 254175
rect 298462 254147 298990 254175
rect -958 254113 298990 254147
rect -958 254085 -430 254113
rect -402 254085 -368 254113
rect -340 254085 -306 254113
rect -278 254085 -244 254113
rect -216 254085 2757 254113
rect 2785 254085 2819 254113
rect 2847 254085 2881 254113
rect 2909 254085 2943 254113
rect 2971 254085 18117 254113
rect 18145 254085 18179 254113
rect 18207 254085 18241 254113
rect 18269 254085 18303 254113
rect 18331 254085 22259 254113
rect 22287 254085 22321 254113
rect 22349 254085 37619 254113
rect 37647 254085 37681 254113
rect 37709 254085 52979 254113
rect 53007 254085 53041 254113
rect 53069 254085 68339 254113
rect 68367 254085 68401 254113
rect 68429 254085 83699 254113
rect 83727 254085 83761 254113
rect 83789 254085 94917 254113
rect 94945 254085 94979 254113
rect 95007 254085 95041 254113
rect 95069 254085 95103 254113
rect 95131 254085 102259 254113
rect 102287 254085 102321 254113
rect 102349 254085 117619 254113
rect 117647 254085 117681 254113
rect 117709 254085 132979 254113
rect 133007 254085 133041 254113
rect 133069 254085 148339 254113
rect 148367 254085 148401 254113
rect 148429 254085 163699 254113
rect 163727 254085 163761 254113
rect 163789 254085 171717 254113
rect 171745 254085 171779 254113
rect 171807 254085 171841 254113
rect 171869 254085 171903 254113
rect 171931 254085 187077 254113
rect 187105 254085 187139 254113
rect 187167 254085 187201 254113
rect 187229 254085 187263 254113
rect 187291 254085 202437 254113
rect 202465 254085 202499 254113
rect 202527 254085 202561 254113
rect 202589 254085 202623 254113
rect 202651 254085 217797 254113
rect 217825 254085 217859 254113
rect 217887 254085 217921 254113
rect 217949 254085 217983 254113
rect 218011 254085 233157 254113
rect 233185 254085 233219 254113
rect 233247 254085 233281 254113
rect 233309 254085 233343 254113
rect 233371 254085 248517 254113
rect 248545 254085 248579 254113
rect 248607 254085 248641 254113
rect 248669 254085 248703 254113
rect 248731 254085 263877 254113
rect 263905 254085 263939 254113
rect 263967 254085 264001 254113
rect 264029 254085 264063 254113
rect 264091 254085 279237 254113
rect 279265 254085 279299 254113
rect 279327 254085 279361 254113
rect 279389 254085 279423 254113
rect 279451 254085 294597 254113
rect 294625 254085 294659 254113
rect 294687 254085 294721 254113
rect 294749 254085 294783 254113
rect 294811 254085 298248 254113
rect 298276 254085 298310 254113
rect 298338 254085 298372 254113
rect 298400 254085 298434 254113
rect 298462 254085 298990 254113
rect -958 254051 298990 254085
rect -958 254023 -430 254051
rect -402 254023 -368 254051
rect -340 254023 -306 254051
rect -278 254023 -244 254051
rect -216 254023 2757 254051
rect 2785 254023 2819 254051
rect 2847 254023 2881 254051
rect 2909 254023 2943 254051
rect 2971 254023 18117 254051
rect 18145 254023 18179 254051
rect 18207 254023 18241 254051
rect 18269 254023 18303 254051
rect 18331 254023 22259 254051
rect 22287 254023 22321 254051
rect 22349 254023 37619 254051
rect 37647 254023 37681 254051
rect 37709 254023 52979 254051
rect 53007 254023 53041 254051
rect 53069 254023 68339 254051
rect 68367 254023 68401 254051
rect 68429 254023 83699 254051
rect 83727 254023 83761 254051
rect 83789 254023 94917 254051
rect 94945 254023 94979 254051
rect 95007 254023 95041 254051
rect 95069 254023 95103 254051
rect 95131 254023 102259 254051
rect 102287 254023 102321 254051
rect 102349 254023 117619 254051
rect 117647 254023 117681 254051
rect 117709 254023 132979 254051
rect 133007 254023 133041 254051
rect 133069 254023 148339 254051
rect 148367 254023 148401 254051
rect 148429 254023 163699 254051
rect 163727 254023 163761 254051
rect 163789 254023 171717 254051
rect 171745 254023 171779 254051
rect 171807 254023 171841 254051
rect 171869 254023 171903 254051
rect 171931 254023 187077 254051
rect 187105 254023 187139 254051
rect 187167 254023 187201 254051
rect 187229 254023 187263 254051
rect 187291 254023 202437 254051
rect 202465 254023 202499 254051
rect 202527 254023 202561 254051
rect 202589 254023 202623 254051
rect 202651 254023 217797 254051
rect 217825 254023 217859 254051
rect 217887 254023 217921 254051
rect 217949 254023 217983 254051
rect 218011 254023 233157 254051
rect 233185 254023 233219 254051
rect 233247 254023 233281 254051
rect 233309 254023 233343 254051
rect 233371 254023 248517 254051
rect 248545 254023 248579 254051
rect 248607 254023 248641 254051
rect 248669 254023 248703 254051
rect 248731 254023 263877 254051
rect 263905 254023 263939 254051
rect 263967 254023 264001 254051
rect 264029 254023 264063 254051
rect 264091 254023 279237 254051
rect 279265 254023 279299 254051
rect 279327 254023 279361 254051
rect 279389 254023 279423 254051
rect 279451 254023 294597 254051
rect 294625 254023 294659 254051
rect 294687 254023 294721 254051
rect 294749 254023 294783 254051
rect 294811 254023 298248 254051
rect 298276 254023 298310 254051
rect 298338 254023 298372 254051
rect 298400 254023 298434 254051
rect 298462 254023 298990 254051
rect -958 253989 298990 254023
rect -958 253961 -430 253989
rect -402 253961 -368 253989
rect -340 253961 -306 253989
rect -278 253961 -244 253989
rect -216 253961 2757 253989
rect 2785 253961 2819 253989
rect 2847 253961 2881 253989
rect 2909 253961 2943 253989
rect 2971 253961 18117 253989
rect 18145 253961 18179 253989
rect 18207 253961 18241 253989
rect 18269 253961 18303 253989
rect 18331 253961 22259 253989
rect 22287 253961 22321 253989
rect 22349 253961 37619 253989
rect 37647 253961 37681 253989
rect 37709 253961 52979 253989
rect 53007 253961 53041 253989
rect 53069 253961 68339 253989
rect 68367 253961 68401 253989
rect 68429 253961 83699 253989
rect 83727 253961 83761 253989
rect 83789 253961 94917 253989
rect 94945 253961 94979 253989
rect 95007 253961 95041 253989
rect 95069 253961 95103 253989
rect 95131 253961 102259 253989
rect 102287 253961 102321 253989
rect 102349 253961 117619 253989
rect 117647 253961 117681 253989
rect 117709 253961 132979 253989
rect 133007 253961 133041 253989
rect 133069 253961 148339 253989
rect 148367 253961 148401 253989
rect 148429 253961 163699 253989
rect 163727 253961 163761 253989
rect 163789 253961 171717 253989
rect 171745 253961 171779 253989
rect 171807 253961 171841 253989
rect 171869 253961 171903 253989
rect 171931 253961 187077 253989
rect 187105 253961 187139 253989
rect 187167 253961 187201 253989
rect 187229 253961 187263 253989
rect 187291 253961 202437 253989
rect 202465 253961 202499 253989
rect 202527 253961 202561 253989
rect 202589 253961 202623 253989
rect 202651 253961 217797 253989
rect 217825 253961 217859 253989
rect 217887 253961 217921 253989
rect 217949 253961 217983 253989
rect 218011 253961 233157 253989
rect 233185 253961 233219 253989
rect 233247 253961 233281 253989
rect 233309 253961 233343 253989
rect 233371 253961 248517 253989
rect 248545 253961 248579 253989
rect 248607 253961 248641 253989
rect 248669 253961 248703 253989
rect 248731 253961 263877 253989
rect 263905 253961 263939 253989
rect 263967 253961 264001 253989
rect 264029 253961 264063 253989
rect 264091 253961 279237 253989
rect 279265 253961 279299 253989
rect 279327 253961 279361 253989
rect 279389 253961 279423 253989
rect 279451 253961 294597 253989
rect 294625 253961 294659 253989
rect 294687 253961 294721 253989
rect 294749 253961 294783 253989
rect 294811 253961 298248 253989
rect 298276 253961 298310 253989
rect 298338 253961 298372 253989
rect 298400 253961 298434 253989
rect 298462 253961 298990 253989
rect -958 253913 298990 253961
rect -958 248175 298990 248223
rect -958 248147 -910 248175
rect -882 248147 -848 248175
rect -820 248147 -786 248175
rect -758 248147 -724 248175
rect -696 248147 4617 248175
rect 4645 248147 4679 248175
rect 4707 248147 4741 248175
rect 4769 248147 4803 248175
rect 4831 248147 29939 248175
rect 29967 248147 30001 248175
rect 30029 248147 45299 248175
rect 45327 248147 45361 248175
rect 45389 248147 60659 248175
rect 60687 248147 60721 248175
rect 60749 248147 76019 248175
rect 76047 248147 76081 248175
rect 76109 248147 96777 248175
rect 96805 248147 96839 248175
rect 96867 248147 96901 248175
rect 96929 248147 96963 248175
rect 96991 248147 109939 248175
rect 109967 248147 110001 248175
rect 110029 248147 125299 248175
rect 125327 248147 125361 248175
rect 125389 248147 140659 248175
rect 140687 248147 140721 248175
rect 140749 248147 156019 248175
rect 156047 248147 156081 248175
rect 156109 248147 173577 248175
rect 173605 248147 173639 248175
rect 173667 248147 173701 248175
rect 173729 248147 173763 248175
rect 173791 248147 188937 248175
rect 188965 248147 188999 248175
rect 189027 248147 189061 248175
rect 189089 248147 189123 248175
rect 189151 248147 204297 248175
rect 204325 248147 204359 248175
rect 204387 248147 204421 248175
rect 204449 248147 204483 248175
rect 204511 248147 219657 248175
rect 219685 248147 219719 248175
rect 219747 248147 219781 248175
rect 219809 248147 219843 248175
rect 219871 248147 235017 248175
rect 235045 248147 235079 248175
rect 235107 248147 235141 248175
rect 235169 248147 235203 248175
rect 235231 248147 250377 248175
rect 250405 248147 250439 248175
rect 250467 248147 250501 248175
rect 250529 248147 250563 248175
rect 250591 248147 265737 248175
rect 265765 248147 265799 248175
rect 265827 248147 265861 248175
rect 265889 248147 265923 248175
rect 265951 248147 281097 248175
rect 281125 248147 281159 248175
rect 281187 248147 281221 248175
rect 281249 248147 281283 248175
rect 281311 248147 296457 248175
rect 296485 248147 296519 248175
rect 296547 248147 296581 248175
rect 296609 248147 296643 248175
rect 296671 248147 298728 248175
rect 298756 248147 298790 248175
rect 298818 248147 298852 248175
rect 298880 248147 298914 248175
rect 298942 248147 298990 248175
rect -958 248113 298990 248147
rect -958 248085 -910 248113
rect -882 248085 -848 248113
rect -820 248085 -786 248113
rect -758 248085 -724 248113
rect -696 248085 4617 248113
rect 4645 248085 4679 248113
rect 4707 248085 4741 248113
rect 4769 248085 4803 248113
rect 4831 248085 29939 248113
rect 29967 248085 30001 248113
rect 30029 248085 45299 248113
rect 45327 248085 45361 248113
rect 45389 248085 60659 248113
rect 60687 248085 60721 248113
rect 60749 248085 76019 248113
rect 76047 248085 76081 248113
rect 76109 248085 96777 248113
rect 96805 248085 96839 248113
rect 96867 248085 96901 248113
rect 96929 248085 96963 248113
rect 96991 248085 109939 248113
rect 109967 248085 110001 248113
rect 110029 248085 125299 248113
rect 125327 248085 125361 248113
rect 125389 248085 140659 248113
rect 140687 248085 140721 248113
rect 140749 248085 156019 248113
rect 156047 248085 156081 248113
rect 156109 248085 173577 248113
rect 173605 248085 173639 248113
rect 173667 248085 173701 248113
rect 173729 248085 173763 248113
rect 173791 248085 188937 248113
rect 188965 248085 188999 248113
rect 189027 248085 189061 248113
rect 189089 248085 189123 248113
rect 189151 248085 204297 248113
rect 204325 248085 204359 248113
rect 204387 248085 204421 248113
rect 204449 248085 204483 248113
rect 204511 248085 219657 248113
rect 219685 248085 219719 248113
rect 219747 248085 219781 248113
rect 219809 248085 219843 248113
rect 219871 248085 235017 248113
rect 235045 248085 235079 248113
rect 235107 248085 235141 248113
rect 235169 248085 235203 248113
rect 235231 248085 250377 248113
rect 250405 248085 250439 248113
rect 250467 248085 250501 248113
rect 250529 248085 250563 248113
rect 250591 248085 265737 248113
rect 265765 248085 265799 248113
rect 265827 248085 265861 248113
rect 265889 248085 265923 248113
rect 265951 248085 281097 248113
rect 281125 248085 281159 248113
rect 281187 248085 281221 248113
rect 281249 248085 281283 248113
rect 281311 248085 296457 248113
rect 296485 248085 296519 248113
rect 296547 248085 296581 248113
rect 296609 248085 296643 248113
rect 296671 248085 298728 248113
rect 298756 248085 298790 248113
rect 298818 248085 298852 248113
rect 298880 248085 298914 248113
rect 298942 248085 298990 248113
rect -958 248051 298990 248085
rect -958 248023 -910 248051
rect -882 248023 -848 248051
rect -820 248023 -786 248051
rect -758 248023 -724 248051
rect -696 248023 4617 248051
rect 4645 248023 4679 248051
rect 4707 248023 4741 248051
rect 4769 248023 4803 248051
rect 4831 248023 29939 248051
rect 29967 248023 30001 248051
rect 30029 248023 45299 248051
rect 45327 248023 45361 248051
rect 45389 248023 60659 248051
rect 60687 248023 60721 248051
rect 60749 248023 76019 248051
rect 76047 248023 76081 248051
rect 76109 248023 96777 248051
rect 96805 248023 96839 248051
rect 96867 248023 96901 248051
rect 96929 248023 96963 248051
rect 96991 248023 109939 248051
rect 109967 248023 110001 248051
rect 110029 248023 125299 248051
rect 125327 248023 125361 248051
rect 125389 248023 140659 248051
rect 140687 248023 140721 248051
rect 140749 248023 156019 248051
rect 156047 248023 156081 248051
rect 156109 248023 173577 248051
rect 173605 248023 173639 248051
rect 173667 248023 173701 248051
rect 173729 248023 173763 248051
rect 173791 248023 188937 248051
rect 188965 248023 188999 248051
rect 189027 248023 189061 248051
rect 189089 248023 189123 248051
rect 189151 248023 204297 248051
rect 204325 248023 204359 248051
rect 204387 248023 204421 248051
rect 204449 248023 204483 248051
rect 204511 248023 219657 248051
rect 219685 248023 219719 248051
rect 219747 248023 219781 248051
rect 219809 248023 219843 248051
rect 219871 248023 235017 248051
rect 235045 248023 235079 248051
rect 235107 248023 235141 248051
rect 235169 248023 235203 248051
rect 235231 248023 250377 248051
rect 250405 248023 250439 248051
rect 250467 248023 250501 248051
rect 250529 248023 250563 248051
rect 250591 248023 265737 248051
rect 265765 248023 265799 248051
rect 265827 248023 265861 248051
rect 265889 248023 265923 248051
rect 265951 248023 281097 248051
rect 281125 248023 281159 248051
rect 281187 248023 281221 248051
rect 281249 248023 281283 248051
rect 281311 248023 296457 248051
rect 296485 248023 296519 248051
rect 296547 248023 296581 248051
rect 296609 248023 296643 248051
rect 296671 248023 298728 248051
rect 298756 248023 298790 248051
rect 298818 248023 298852 248051
rect 298880 248023 298914 248051
rect 298942 248023 298990 248051
rect -958 247989 298990 248023
rect -958 247961 -910 247989
rect -882 247961 -848 247989
rect -820 247961 -786 247989
rect -758 247961 -724 247989
rect -696 247961 4617 247989
rect 4645 247961 4679 247989
rect 4707 247961 4741 247989
rect 4769 247961 4803 247989
rect 4831 247961 29939 247989
rect 29967 247961 30001 247989
rect 30029 247961 45299 247989
rect 45327 247961 45361 247989
rect 45389 247961 60659 247989
rect 60687 247961 60721 247989
rect 60749 247961 76019 247989
rect 76047 247961 76081 247989
rect 76109 247961 96777 247989
rect 96805 247961 96839 247989
rect 96867 247961 96901 247989
rect 96929 247961 96963 247989
rect 96991 247961 109939 247989
rect 109967 247961 110001 247989
rect 110029 247961 125299 247989
rect 125327 247961 125361 247989
rect 125389 247961 140659 247989
rect 140687 247961 140721 247989
rect 140749 247961 156019 247989
rect 156047 247961 156081 247989
rect 156109 247961 173577 247989
rect 173605 247961 173639 247989
rect 173667 247961 173701 247989
rect 173729 247961 173763 247989
rect 173791 247961 188937 247989
rect 188965 247961 188999 247989
rect 189027 247961 189061 247989
rect 189089 247961 189123 247989
rect 189151 247961 204297 247989
rect 204325 247961 204359 247989
rect 204387 247961 204421 247989
rect 204449 247961 204483 247989
rect 204511 247961 219657 247989
rect 219685 247961 219719 247989
rect 219747 247961 219781 247989
rect 219809 247961 219843 247989
rect 219871 247961 235017 247989
rect 235045 247961 235079 247989
rect 235107 247961 235141 247989
rect 235169 247961 235203 247989
rect 235231 247961 250377 247989
rect 250405 247961 250439 247989
rect 250467 247961 250501 247989
rect 250529 247961 250563 247989
rect 250591 247961 265737 247989
rect 265765 247961 265799 247989
rect 265827 247961 265861 247989
rect 265889 247961 265923 247989
rect 265951 247961 281097 247989
rect 281125 247961 281159 247989
rect 281187 247961 281221 247989
rect 281249 247961 281283 247989
rect 281311 247961 296457 247989
rect 296485 247961 296519 247989
rect 296547 247961 296581 247989
rect 296609 247961 296643 247989
rect 296671 247961 298728 247989
rect 298756 247961 298790 247989
rect 298818 247961 298852 247989
rect 298880 247961 298914 247989
rect 298942 247961 298990 247989
rect -958 247913 298990 247961
rect -958 245175 298990 245223
rect -958 245147 -430 245175
rect -402 245147 -368 245175
rect -340 245147 -306 245175
rect -278 245147 -244 245175
rect -216 245147 2757 245175
rect 2785 245147 2819 245175
rect 2847 245147 2881 245175
rect 2909 245147 2943 245175
rect 2971 245147 18117 245175
rect 18145 245147 18179 245175
rect 18207 245147 18241 245175
rect 18269 245147 18303 245175
rect 18331 245147 22259 245175
rect 22287 245147 22321 245175
rect 22349 245147 37619 245175
rect 37647 245147 37681 245175
rect 37709 245147 52979 245175
rect 53007 245147 53041 245175
rect 53069 245147 68339 245175
rect 68367 245147 68401 245175
rect 68429 245147 83699 245175
rect 83727 245147 83761 245175
rect 83789 245147 94917 245175
rect 94945 245147 94979 245175
rect 95007 245147 95041 245175
rect 95069 245147 95103 245175
rect 95131 245147 102259 245175
rect 102287 245147 102321 245175
rect 102349 245147 117619 245175
rect 117647 245147 117681 245175
rect 117709 245147 132979 245175
rect 133007 245147 133041 245175
rect 133069 245147 148339 245175
rect 148367 245147 148401 245175
rect 148429 245147 163699 245175
rect 163727 245147 163761 245175
rect 163789 245147 171717 245175
rect 171745 245147 171779 245175
rect 171807 245147 171841 245175
rect 171869 245147 171903 245175
rect 171931 245147 187077 245175
rect 187105 245147 187139 245175
rect 187167 245147 187201 245175
rect 187229 245147 187263 245175
rect 187291 245147 202437 245175
rect 202465 245147 202499 245175
rect 202527 245147 202561 245175
rect 202589 245147 202623 245175
rect 202651 245147 217797 245175
rect 217825 245147 217859 245175
rect 217887 245147 217921 245175
rect 217949 245147 217983 245175
rect 218011 245147 233157 245175
rect 233185 245147 233219 245175
rect 233247 245147 233281 245175
rect 233309 245147 233343 245175
rect 233371 245147 248517 245175
rect 248545 245147 248579 245175
rect 248607 245147 248641 245175
rect 248669 245147 248703 245175
rect 248731 245147 263877 245175
rect 263905 245147 263939 245175
rect 263967 245147 264001 245175
rect 264029 245147 264063 245175
rect 264091 245147 279237 245175
rect 279265 245147 279299 245175
rect 279327 245147 279361 245175
rect 279389 245147 279423 245175
rect 279451 245147 294597 245175
rect 294625 245147 294659 245175
rect 294687 245147 294721 245175
rect 294749 245147 294783 245175
rect 294811 245147 298248 245175
rect 298276 245147 298310 245175
rect 298338 245147 298372 245175
rect 298400 245147 298434 245175
rect 298462 245147 298990 245175
rect -958 245113 298990 245147
rect -958 245085 -430 245113
rect -402 245085 -368 245113
rect -340 245085 -306 245113
rect -278 245085 -244 245113
rect -216 245085 2757 245113
rect 2785 245085 2819 245113
rect 2847 245085 2881 245113
rect 2909 245085 2943 245113
rect 2971 245085 18117 245113
rect 18145 245085 18179 245113
rect 18207 245085 18241 245113
rect 18269 245085 18303 245113
rect 18331 245085 22259 245113
rect 22287 245085 22321 245113
rect 22349 245085 37619 245113
rect 37647 245085 37681 245113
rect 37709 245085 52979 245113
rect 53007 245085 53041 245113
rect 53069 245085 68339 245113
rect 68367 245085 68401 245113
rect 68429 245085 83699 245113
rect 83727 245085 83761 245113
rect 83789 245085 94917 245113
rect 94945 245085 94979 245113
rect 95007 245085 95041 245113
rect 95069 245085 95103 245113
rect 95131 245085 102259 245113
rect 102287 245085 102321 245113
rect 102349 245085 117619 245113
rect 117647 245085 117681 245113
rect 117709 245085 132979 245113
rect 133007 245085 133041 245113
rect 133069 245085 148339 245113
rect 148367 245085 148401 245113
rect 148429 245085 163699 245113
rect 163727 245085 163761 245113
rect 163789 245085 171717 245113
rect 171745 245085 171779 245113
rect 171807 245085 171841 245113
rect 171869 245085 171903 245113
rect 171931 245085 187077 245113
rect 187105 245085 187139 245113
rect 187167 245085 187201 245113
rect 187229 245085 187263 245113
rect 187291 245085 202437 245113
rect 202465 245085 202499 245113
rect 202527 245085 202561 245113
rect 202589 245085 202623 245113
rect 202651 245085 217797 245113
rect 217825 245085 217859 245113
rect 217887 245085 217921 245113
rect 217949 245085 217983 245113
rect 218011 245085 233157 245113
rect 233185 245085 233219 245113
rect 233247 245085 233281 245113
rect 233309 245085 233343 245113
rect 233371 245085 248517 245113
rect 248545 245085 248579 245113
rect 248607 245085 248641 245113
rect 248669 245085 248703 245113
rect 248731 245085 263877 245113
rect 263905 245085 263939 245113
rect 263967 245085 264001 245113
rect 264029 245085 264063 245113
rect 264091 245085 279237 245113
rect 279265 245085 279299 245113
rect 279327 245085 279361 245113
rect 279389 245085 279423 245113
rect 279451 245085 294597 245113
rect 294625 245085 294659 245113
rect 294687 245085 294721 245113
rect 294749 245085 294783 245113
rect 294811 245085 298248 245113
rect 298276 245085 298310 245113
rect 298338 245085 298372 245113
rect 298400 245085 298434 245113
rect 298462 245085 298990 245113
rect -958 245051 298990 245085
rect -958 245023 -430 245051
rect -402 245023 -368 245051
rect -340 245023 -306 245051
rect -278 245023 -244 245051
rect -216 245023 2757 245051
rect 2785 245023 2819 245051
rect 2847 245023 2881 245051
rect 2909 245023 2943 245051
rect 2971 245023 18117 245051
rect 18145 245023 18179 245051
rect 18207 245023 18241 245051
rect 18269 245023 18303 245051
rect 18331 245023 22259 245051
rect 22287 245023 22321 245051
rect 22349 245023 37619 245051
rect 37647 245023 37681 245051
rect 37709 245023 52979 245051
rect 53007 245023 53041 245051
rect 53069 245023 68339 245051
rect 68367 245023 68401 245051
rect 68429 245023 83699 245051
rect 83727 245023 83761 245051
rect 83789 245023 94917 245051
rect 94945 245023 94979 245051
rect 95007 245023 95041 245051
rect 95069 245023 95103 245051
rect 95131 245023 102259 245051
rect 102287 245023 102321 245051
rect 102349 245023 117619 245051
rect 117647 245023 117681 245051
rect 117709 245023 132979 245051
rect 133007 245023 133041 245051
rect 133069 245023 148339 245051
rect 148367 245023 148401 245051
rect 148429 245023 163699 245051
rect 163727 245023 163761 245051
rect 163789 245023 171717 245051
rect 171745 245023 171779 245051
rect 171807 245023 171841 245051
rect 171869 245023 171903 245051
rect 171931 245023 187077 245051
rect 187105 245023 187139 245051
rect 187167 245023 187201 245051
rect 187229 245023 187263 245051
rect 187291 245023 202437 245051
rect 202465 245023 202499 245051
rect 202527 245023 202561 245051
rect 202589 245023 202623 245051
rect 202651 245023 217797 245051
rect 217825 245023 217859 245051
rect 217887 245023 217921 245051
rect 217949 245023 217983 245051
rect 218011 245023 233157 245051
rect 233185 245023 233219 245051
rect 233247 245023 233281 245051
rect 233309 245023 233343 245051
rect 233371 245023 248517 245051
rect 248545 245023 248579 245051
rect 248607 245023 248641 245051
rect 248669 245023 248703 245051
rect 248731 245023 263877 245051
rect 263905 245023 263939 245051
rect 263967 245023 264001 245051
rect 264029 245023 264063 245051
rect 264091 245023 279237 245051
rect 279265 245023 279299 245051
rect 279327 245023 279361 245051
rect 279389 245023 279423 245051
rect 279451 245023 294597 245051
rect 294625 245023 294659 245051
rect 294687 245023 294721 245051
rect 294749 245023 294783 245051
rect 294811 245023 298248 245051
rect 298276 245023 298310 245051
rect 298338 245023 298372 245051
rect 298400 245023 298434 245051
rect 298462 245023 298990 245051
rect -958 244989 298990 245023
rect -958 244961 -430 244989
rect -402 244961 -368 244989
rect -340 244961 -306 244989
rect -278 244961 -244 244989
rect -216 244961 2757 244989
rect 2785 244961 2819 244989
rect 2847 244961 2881 244989
rect 2909 244961 2943 244989
rect 2971 244961 18117 244989
rect 18145 244961 18179 244989
rect 18207 244961 18241 244989
rect 18269 244961 18303 244989
rect 18331 244961 22259 244989
rect 22287 244961 22321 244989
rect 22349 244961 37619 244989
rect 37647 244961 37681 244989
rect 37709 244961 52979 244989
rect 53007 244961 53041 244989
rect 53069 244961 68339 244989
rect 68367 244961 68401 244989
rect 68429 244961 83699 244989
rect 83727 244961 83761 244989
rect 83789 244961 94917 244989
rect 94945 244961 94979 244989
rect 95007 244961 95041 244989
rect 95069 244961 95103 244989
rect 95131 244961 102259 244989
rect 102287 244961 102321 244989
rect 102349 244961 117619 244989
rect 117647 244961 117681 244989
rect 117709 244961 132979 244989
rect 133007 244961 133041 244989
rect 133069 244961 148339 244989
rect 148367 244961 148401 244989
rect 148429 244961 163699 244989
rect 163727 244961 163761 244989
rect 163789 244961 171717 244989
rect 171745 244961 171779 244989
rect 171807 244961 171841 244989
rect 171869 244961 171903 244989
rect 171931 244961 187077 244989
rect 187105 244961 187139 244989
rect 187167 244961 187201 244989
rect 187229 244961 187263 244989
rect 187291 244961 202437 244989
rect 202465 244961 202499 244989
rect 202527 244961 202561 244989
rect 202589 244961 202623 244989
rect 202651 244961 217797 244989
rect 217825 244961 217859 244989
rect 217887 244961 217921 244989
rect 217949 244961 217983 244989
rect 218011 244961 233157 244989
rect 233185 244961 233219 244989
rect 233247 244961 233281 244989
rect 233309 244961 233343 244989
rect 233371 244961 248517 244989
rect 248545 244961 248579 244989
rect 248607 244961 248641 244989
rect 248669 244961 248703 244989
rect 248731 244961 263877 244989
rect 263905 244961 263939 244989
rect 263967 244961 264001 244989
rect 264029 244961 264063 244989
rect 264091 244961 279237 244989
rect 279265 244961 279299 244989
rect 279327 244961 279361 244989
rect 279389 244961 279423 244989
rect 279451 244961 294597 244989
rect 294625 244961 294659 244989
rect 294687 244961 294721 244989
rect 294749 244961 294783 244989
rect 294811 244961 298248 244989
rect 298276 244961 298310 244989
rect 298338 244961 298372 244989
rect 298400 244961 298434 244989
rect 298462 244961 298990 244989
rect -958 244913 298990 244961
rect -958 239175 298990 239223
rect -958 239147 -910 239175
rect -882 239147 -848 239175
rect -820 239147 -786 239175
rect -758 239147 -724 239175
rect -696 239147 4617 239175
rect 4645 239147 4679 239175
rect 4707 239147 4741 239175
rect 4769 239147 4803 239175
rect 4831 239147 29939 239175
rect 29967 239147 30001 239175
rect 30029 239147 45299 239175
rect 45327 239147 45361 239175
rect 45389 239147 60659 239175
rect 60687 239147 60721 239175
rect 60749 239147 76019 239175
rect 76047 239147 76081 239175
rect 76109 239147 96777 239175
rect 96805 239147 96839 239175
rect 96867 239147 96901 239175
rect 96929 239147 96963 239175
rect 96991 239147 109939 239175
rect 109967 239147 110001 239175
rect 110029 239147 125299 239175
rect 125327 239147 125361 239175
rect 125389 239147 140659 239175
rect 140687 239147 140721 239175
rect 140749 239147 156019 239175
rect 156047 239147 156081 239175
rect 156109 239147 173577 239175
rect 173605 239147 173639 239175
rect 173667 239147 173701 239175
rect 173729 239147 173763 239175
rect 173791 239147 188937 239175
rect 188965 239147 188999 239175
rect 189027 239147 189061 239175
rect 189089 239147 189123 239175
rect 189151 239147 204297 239175
rect 204325 239147 204359 239175
rect 204387 239147 204421 239175
rect 204449 239147 204483 239175
rect 204511 239147 219657 239175
rect 219685 239147 219719 239175
rect 219747 239147 219781 239175
rect 219809 239147 219843 239175
rect 219871 239147 235017 239175
rect 235045 239147 235079 239175
rect 235107 239147 235141 239175
rect 235169 239147 235203 239175
rect 235231 239147 250377 239175
rect 250405 239147 250439 239175
rect 250467 239147 250501 239175
rect 250529 239147 250563 239175
rect 250591 239147 265737 239175
rect 265765 239147 265799 239175
rect 265827 239147 265861 239175
rect 265889 239147 265923 239175
rect 265951 239147 281097 239175
rect 281125 239147 281159 239175
rect 281187 239147 281221 239175
rect 281249 239147 281283 239175
rect 281311 239147 296457 239175
rect 296485 239147 296519 239175
rect 296547 239147 296581 239175
rect 296609 239147 296643 239175
rect 296671 239147 298728 239175
rect 298756 239147 298790 239175
rect 298818 239147 298852 239175
rect 298880 239147 298914 239175
rect 298942 239147 298990 239175
rect -958 239113 298990 239147
rect -958 239085 -910 239113
rect -882 239085 -848 239113
rect -820 239085 -786 239113
rect -758 239085 -724 239113
rect -696 239085 4617 239113
rect 4645 239085 4679 239113
rect 4707 239085 4741 239113
rect 4769 239085 4803 239113
rect 4831 239085 29939 239113
rect 29967 239085 30001 239113
rect 30029 239085 45299 239113
rect 45327 239085 45361 239113
rect 45389 239085 60659 239113
rect 60687 239085 60721 239113
rect 60749 239085 76019 239113
rect 76047 239085 76081 239113
rect 76109 239085 96777 239113
rect 96805 239085 96839 239113
rect 96867 239085 96901 239113
rect 96929 239085 96963 239113
rect 96991 239085 109939 239113
rect 109967 239085 110001 239113
rect 110029 239085 125299 239113
rect 125327 239085 125361 239113
rect 125389 239085 140659 239113
rect 140687 239085 140721 239113
rect 140749 239085 156019 239113
rect 156047 239085 156081 239113
rect 156109 239085 173577 239113
rect 173605 239085 173639 239113
rect 173667 239085 173701 239113
rect 173729 239085 173763 239113
rect 173791 239085 188937 239113
rect 188965 239085 188999 239113
rect 189027 239085 189061 239113
rect 189089 239085 189123 239113
rect 189151 239085 204297 239113
rect 204325 239085 204359 239113
rect 204387 239085 204421 239113
rect 204449 239085 204483 239113
rect 204511 239085 219657 239113
rect 219685 239085 219719 239113
rect 219747 239085 219781 239113
rect 219809 239085 219843 239113
rect 219871 239085 235017 239113
rect 235045 239085 235079 239113
rect 235107 239085 235141 239113
rect 235169 239085 235203 239113
rect 235231 239085 250377 239113
rect 250405 239085 250439 239113
rect 250467 239085 250501 239113
rect 250529 239085 250563 239113
rect 250591 239085 265737 239113
rect 265765 239085 265799 239113
rect 265827 239085 265861 239113
rect 265889 239085 265923 239113
rect 265951 239085 281097 239113
rect 281125 239085 281159 239113
rect 281187 239085 281221 239113
rect 281249 239085 281283 239113
rect 281311 239085 296457 239113
rect 296485 239085 296519 239113
rect 296547 239085 296581 239113
rect 296609 239085 296643 239113
rect 296671 239085 298728 239113
rect 298756 239085 298790 239113
rect 298818 239085 298852 239113
rect 298880 239085 298914 239113
rect 298942 239085 298990 239113
rect -958 239051 298990 239085
rect -958 239023 -910 239051
rect -882 239023 -848 239051
rect -820 239023 -786 239051
rect -758 239023 -724 239051
rect -696 239023 4617 239051
rect 4645 239023 4679 239051
rect 4707 239023 4741 239051
rect 4769 239023 4803 239051
rect 4831 239023 29939 239051
rect 29967 239023 30001 239051
rect 30029 239023 45299 239051
rect 45327 239023 45361 239051
rect 45389 239023 60659 239051
rect 60687 239023 60721 239051
rect 60749 239023 76019 239051
rect 76047 239023 76081 239051
rect 76109 239023 96777 239051
rect 96805 239023 96839 239051
rect 96867 239023 96901 239051
rect 96929 239023 96963 239051
rect 96991 239023 109939 239051
rect 109967 239023 110001 239051
rect 110029 239023 125299 239051
rect 125327 239023 125361 239051
rect 125389 239023 140659 239051
rect 140687 239023 140721 239051
rect 140749 239023 156019 239051
rect 156047 239023 156081 239051
rect 156109 239023 173577 239051
rect 173605 239023 173639 239051
rect 173667 239023 173701 239051
rect 173729 239023 173763 239051
rect 173791 239023 188937 239051
rect 188965 239023 188999 239051
rect 189027 239023 189061 239051
rect 189089 239023 189123 239051
rect 189151 239023 204297 239051
rect 204325 239023 204359 239051
rect 204387 239023 204421 239051
rect 204449 239023 204483 239051
rect 204511 239023 219657 239051
rect 219685 239023 219719 239051
rect 219747 239023 219781 239051
rect 219809 239023 219843 239051
rect 219871 239023 235017 239051
rect 235045 239023 235079 239051
rect 235107 239023 235141 239051
rect 235169 239023 235203 239051
rect 235231 239023 250377 239051
rect 250405 239023 250439 239051
rect 250467 239023 250501 239051
rect 250529 239023 250563 239051
rect 250591 239023 265737 239051
rect 265765 239023 265799 239051
rect 265827 239023 265861 239051
rect 265889 239023 265923 239051
rect 265951 239023 281097 239051
rect 281125 239023 281159 239051
rect 281187 239023 281221 239051
rect 281249 239023 281283 239051
rect 281311 239023 296457 239051
rect 296485 239023 296519 239051
rect 296547 239023 296581 239051
rect 296609 239023 296643 239051
rect 296671 239023 298728 239051
rect 298756 239023 298790 239051
rect 298818 239023 298852 239051
rect 298880 239023 298914 239051
rect 298942 239023 298990 239051
rect -958 238989 298990 239023
rect -958 238961 -910 238989
rect -882 238961 -848 238989
rect -820 238961 -786 238989
rect -758 238961 -724 238989
rect -696 238961 4617 238989
rect 4645 238961 4679 238989
rect 4707 238961 4741 238989
rect 4769 238961 4803 238989
rect 4831 238961 29939 238989
rect 29967 238961 30001 238989
rect 30029 238961 45299 238989
rect 45327 238961 45361 238989
rect 45389 238961 60659 238989
rect 60687 238961 60721 238989
rect 60749 238961 76019 238989
rect 76047 238961 76081 238989
rect 76109 238961 96777 238989
rect 96805 238961 96839 238989
rect 96867 238961 96901 238989
rect 96929 238961 96963 238989
rect 96991 238961 109939 238989
rect 109967 238961 110001 238989
rect 110029 238961 125299 238989
rect 125327 238961 125361 238989
rect 125389 238961 140659 238989
rect 140687 238961 140721 238989
rect 140749 238961 156019 238989
rect 156047 238961 156081 238989
rect 156109 238961 173577 238989
rect 173605 238961 173639 238989
rect 173667 238961 173701 238989
rect 173729 238961 173763 238989
rect 173791 238961 188937 238989
rect 188965 238961 188999 238989
rect 189027 238961 189061 238989
rect 189089 238961 189123 238989
rect 189151 238961 204297 238989
rect 204325 238961 204359 238989
rect 204387 238961 204421 238989
rect 204449 238961 204483 238989
rect 204511 238961 219657 238989
rect 219685 238961 219719 238989
rect 219747 238961 219781 238989
rect 219809 238961 219843 238989
rect 219871 238961 235017 238989
rect 235045 238961 235079 238989
rect 235107 238961 235141 238989
rect 235169 238961 235203 238989
rect 235231 238961 250377 238989
rect 250405 238961 250439 238989
rect 250467 238961 250501 238989
rect 250529 238961 250563 238989
rect 250591 238961 265737 238989
rect 265765 238961 265799 238989
rect 265827 238961 265861 238989
rect 265889 238961 265923 238989
rect 265951 238961 281097 238989
rect 281125 238961 281159 238989
rect 281187 238961 281221 238989
rect 281249 238961 281283 238989
rect 281311 238961 296457 238989
rect 296485 238961 296519 238989
rect 296547 238961 296581 238989
rect 296609 238961 296643 238989
rect 296671 238961 298728 238989
rect 298756 238961 298790 238989
rect 298818 238961 298852 238989
rect 298880 238961 298914 238989
rect 298942 238961 298990 238989
rect -958 238913 298990 238961
rect -958 236175 298990 236223
rect -958 236147 -430 236175
rect -402 236147 -368 236175
rect -340 236147 -306 236175
rect -278 236147 -244 236175
rect -216 236147 2757 236175
rect 2785 236147 2819 236175
rect 2847 236147 2881 236175
rect 2909 236147 2943 236175
rect 2971 236147 18117 236175
rect 18145 236147 18179 236175
rect 18207 236147 18241 236175
rect 18269 236147 18303 236175
rect 18331 236147 22259 236175
rect 22287 236147 22321 236175
rect 22349 236147 37619 236175
rect 37647 236147 37681 236175
rect 37709 236147 52979 236175
rect 53007 236147 53041 236175
rect 53069 236147 68339 236175
rect 68367 236147 68401 236175
rect 68429 236147 83699 236175
rect 83727 236147 83761 236175
rect 83789 236147 94917 236175
rect 94945 236147 94979 236175
rect 95007 236147 95041 236175
rect 95069 236147 95103 236175
rect 95131 236147 102259 236175
rect 102287 236147 102321 236175
rect 102349 236147 117619 236175
rect 117647 236147 117681 236175
rect 117709 236147 132979 236175
rect 133007 236147 133041 236175
rect 133069 236147 148339 236175
rect 148367 236147 148401 236175
rect 148429 236147 163699 236175
rect 163727 236147 163761 236175
rect 163789 236147 171717 236175
rect 171745 236147 171779 236175
rect 171807 236147 171841 236175
rect 171869 236147 171903 236175
rect 171931 236147 187077 236175
rect 187105 236147 187139 236175
rect 187167 236147 187201 236175
rect 187229 236147 187263 236175
rect 187291 236147 202437 236175
rect 202465 236147 202499 236175
rect 202527 236147 202561 236175
rect 202589 236147 202623 236175
rect 202651 236147 217797 236175
rect 217825 236147 217859 236175
rect 217887 236147 217921 236175
rect 217949 236147 217983 236175
rect 218011 236147 233157 236175
rect 233185 236147 233219 236175
rect 233247 236147 233281 236175
rect 233309 236147 233343 236175
rect 233371 236147 248517 236175
rect 248545 236147 248579 236175
rect 248607 236147 248641 236175
rect 248669 236147 248703 236175
rect 248731 236147 263877 236175
rect 263905 236147 263939 236175
rect 263967 236147 264001 236175
rect 264029 236147 264063 236175
rect 264091 236147 279237 236175
rect 279265 236147 279299 236175
rect 279327 236147 279361 236175
rect 279389 236147 279423 236175
rect 279451 236147 294597 236175
rect 294625 236147 294659 236175
rect 294687 236147 294721 236175
rect 294749 236147 294783 236175
rect 294811 236147 298248 236175
rect 298276 236147 298310 236175
rect 298338 236147 298372 236175
rect 298400 236147 298434 236175
rect 298462 236147 298990 236175
rect -958 236113 298990 236147
rect -958 236085 -430 236113
rect -402 236085 -368 236113
rect -340 236085 -306 236113
rect -278 236085 -244 236113
rect -216 236085 2757 236113
rect 2785 236085 2819 236113
rect 2847 236085 2881 236113
rect 2909 236085 2943 236113
rect 2971 236085 18117 236113
rect 18145 236085 18179 236113
rect 18207 236085 18241 236113
rect 18269 236085 18303 236113
rect 18331 236085 22259 236113
rect 22287 236085 22321 236113
rect 22349 236085 37619 236113
rect 37647 236085 37681 236113
rect 37709 236085 52979 236113
rect 53007 236085 53041 236113
rect 53069 236085 68339 236113
rect 68367 236085 68401 236113
rect 68429 236085 83699 236113
rect 83727 236085 83761 236113
rect 83789 236085 94917 236113
rect 94945 236085 94979 236113
rect 95007 236085 95041 236113
rect 95069 236085 95103 236113
rect 95131 236085 102259 236113
rect 102287 236085 102321 236113
rect 102349 236085 117619 236113
rect 117647 236085 117681 236113
rect 117709 236085 132979 236113
rect 133007 236085 133041 236113
rect 133069 236085 148339 236113
rect 148367 236085 148401 236113
rect 148429 236085 163699 236113
rect 163727 236085 163761 236113
rect 163789 236085 171717 236113
rect 171745 236085 171779 236113
rect 171807 236085 171841 236113
rect 171869 236085 171903 236113
rect 171931 236085 187077 236113
rect 187105 236085 187139 236113
rect 187167 236085 187201 236113
rect 187229 236085 187263 236113
rect 187291 236085 202437 236113
rect 202465 236085 202499 236113
rect 202527 236085 202561 236113
rect 202589 236085 202623 236113
rect 202651 236085 217797 236113
rect 217825 236085 217859 236113
rect 217887 236085 217921 236113
rect 217949 236085 217983 236113
rect 218011 236085 233157 236113
rect 233185 236085 233219 236113
rect 233247 236085 233281 236113
rect 233309 236085 233343 236113
rect 233371 236085 248517 236113
rect 248545 236085 248579 236113
rect 248607 236085 248641 236113
rect 248669 236085 248703 236113
rect 248731 236085 263877 236113
rect 263905 236085 263939 236113
rect 263967 236085 264001 236113
rect 264029 236085 264063 236113
rect 264091 236085 279237 236113
rect 279265 236085 279299 236113
rect 279327 236085 279361 236113
rect 279389 236085 279423 236113
rect 279451 236085 294597 236113
rect 294625 236085 294659 236113
rect 294687 236085 294721 236113
rect 294749 236085 294783 236113
rect 294811 236085 298248 236113
rect 298276 236085 298310 236113
rect 298338 236085 298372 236113
rect 298400 236085 298434 236113
rect 298462 236085 298990 236113
rect -958 236051 298990 236085
rect -958 236023 -430 236051
rect -402 236023 -368 236051
rect -340 236023 -306 236051
rect -278 236023 -244 236051
rect -216 236023 2757 236051
rect 2785 236023 2819 236051
rect 2847 236023 2881 236051
rect 2909 236023 2943 236051
rect 2971 236023 18117 236051
rect 18145 236023 18179 236051
rect 18207 236023 18241 236051
rect 18269 236023 18303 236051
rect 18331 236023 22259 236051
rect 22287 236023 22321 236051
rect 22349 236023 37619 236051
rect 37647 236023 37681 236051
rect 37709 236023 52979 236051
rect 53007 236023 53041 236051
rect 53069 236023 68339 236051
rect 68367 236023 68401 236051
rect 68429 236023 83699 236051
rect 83727 236023 83761 236051
rect 83789 236023 94917 236051
rect 94945 236023 94979 236051
rect 95007 236023 95041 236051
rect 95069 236023 95103 236051
rect 95131 236023 102259 236051
rect 102287 236023 102321 236051
rect 102349 236023 117619 236051
rect 117647 236023 117681 236051
rect 117709 236023 132979 236051
rect 133007 236023 133041 236051
rect 133069 236023 148339 236051
rect 148367 236023 148401 236051
rect 148429 236023 163699 236051
rect 163727 236023 163761 236051
rect 163789 236023 171717 236051
rect 171745 236023 171779 236051
rect 171807 236023 171841 236051
rect 171869 236023 171903 236051
rect 171931 236023 187077 236051
rect 187105 236023 187139 236051
rect 187167 236023 187201 236051
rect 187229 236023 187263 236051
rect 187291 236023 202437 236051
rect 202465 236023 202499 236051
rect 202527 236023 202561 236051
rect 202589 236023 202623 236051
rect 202651 236023 217797 236051
rect 217825 236023 217859 236051
rect 217887 236023 217921 236051
rect 217949 236023 217983 236051
rect 218011 236023 233157 236051
rect 233185 236023 233219 236051
rect 233247 236023 233281 236051
rect 233309 236023 233343 236051
rect 233371 236023 248517 236051
rect 248545 236023 248579 236051
rect 248607 236023 248641 236051
rect 248669 236023 248703 236051
rect 248731 236023 263877 236051
rect 263905 236023 263939 236051
rect 263967 236023 264001 236051
rect 264029 236023 264063 236051
rect 264091 236023 279237 236051
rect 279265 236023 279299 236051
rect 279327 236023 279361 236051
rect 279389 236023 279423 236051
rect 279451 236023 294597 236051
rect 294625 236023 294659 236051
rect 294687 236023 294721 236051
rect 294749 236023 294783 236051
rect 294811 236023 298248 236051
rect 298276 236023 298310 236051
rect 298338 236023 298372 236051
rect 298400 236023 298434 236051
rect 298462 236023 298990 236051
rect -958 235989 298990 236023
rect -958 235961 -430 235989
rect -402 235961 -368 235989
rect -340 235961 -306 235989
rect -278 235961 -244 235989
rect -216 235961 2757 235989
rect 2785 235961 2819 235989
rect 2847 235961 2881 235989
rect 2909 235961 2943 235989
rect 2971 235961 18117 235989
rect 18145 235961 18179 235989
rect 18207 235961 18241 235989
rect 18269 235961 18303 235989
rect 18331 235961 22259 235989
rect 22287 235961 22321 235989
rect 22349 235961 37619 235989
rect 37647 235961 37681 235989
rect 37709 235961 52979 235989
rect 53007 235961 53041 235989
rect 53069 235961 68339 235989
rect 68367 235961 68401 235989
rect 68429 235961 83699 235989
rect 83727 235961 83761 235989
rect 83789 235961 94917 235989
rect 94945 235961 94979 235989
rect 95007 235961 95041 235989
rect 95069 235961 95103 235989
rect 95131 235961 102259 235989
rect 102287 235961 102321 235989
rect 102349 235961 117619 235989
rect 117647 235961 117681 235989
rect 117709 235961 132979 235989
rect 133007 235961 133041 235989
rect 133069 235961 148339 235989
rect 148367 235961 148401 235989
rect 148429 235961 163699 235989
rect 163727 235961 163761 235989
rect 163789 235961 171717 235989
rect 171745 235961 171779 235989
rect 171807 235961 171841 235989
rect 171869 235961 171903 235989
rect 171931 235961 187077 235989
rect 187105 235961 187139 235989
rect 187167 235961 187201 235989
rect 187229 235961 187263 235989
rect 187291 235961 202437 235989
rect 202465 235961 202499 235989
rect 202527 235961 202561 235989
rect 202589 235961 202623 235989
rect 202651 235961 217797 235989
rect 217825 235961 217859 235989
rect 217887 235961 217921 235989
rect 217949 235961 217983 235989
rect 218011 235961 233157 235989
rect 233185 235961 233219 235989
rect 233247 235961 233281 235989
rect 233309 235961 233343 235989
rect 233371 235961 248517 235989
rect 248545 235961 248579 235989
rect 248607 235961 248641 235989
rect 248669 235961 248703 235989
rect 248731 235961 263877 235989
rect 263905 235961 263939 235989
rect 263967 235961 264001 235989
rect 264029 235961 264063 235989
rect 264091 235961 279237 235989
rect 279265 235961 279299 235989
rect 279327 235961 279361 235989
rect 279389 235961 279423 235989
rect 279451 235961 294597 235989
rect 294625 235961 294659 235989
rect 294687 235961 294721 235989
rect 294749 235961 294783 235989
rect 294811 235961 298248 235989
rect 298276 235961 298310 235989
rect 298338 235961 298372 235989
rect 298400 235961 298434 235989
rect 298462 235961 298990 235989
rect -958 235913 298990 235961
rect -958 230175 298990 230223
rect -958 230147 -910 230175
rect -882 230147 -848 230175
rect -820 230147 -786 230175
rect -758 230147 -724 230175
rect -696 230147 4617 230175
rect 4645 230147 4679 230175
rect 4707 230147 4741 230175
rect 4769 230147 4803 230175
rect 4831 230147 29939 230175
rect 29967 230147 30001 230175
rect 30029 230147 45299 230175
rect 45327 230147 45361 230175
rect 45389 230147 60659 230175
rect 60687 230147 60721 230175
rect 60749 230147 76019 230175
rect 76047 230147 76081 230175
rect 76109 230147 96777 230175
rect 96805 230147 96839 230175
rect 96867 230147 96901 230175
rect 96929 230147 96963 230175
rect 96991 230147 109939 230175
rect 109967 230147 110001 230175
rect 110029 230147 125299 230175
rect 125327 230147 125361 230175
rect 125389 230147 140659 230175
rect 140687 230147 140721 230175
rect 140749 230147 156019 230175
rect 156047 230147 156081 230175
rect 156109 230147 173577 230175
rect 173605 230147 173639 230175
rect 173667 230147 173701 230175
rect 173729 230147 173763 230175
rect 173791 230147 188937 230175
rect 188965 230147 188999 230175
rect 189027 230147 189061 230175
rect 189089 230147 189123 230175
rect 189151 230147 204297 230175
rect 204325 230147 204359 230175
rect 204387 230147 204421 230175
rect 204449 230147 204483 230175
rect 204511 230147 219657 230175
rect 219685 230147 219719 230175
rect 219747 230147 219781 230175
rect 219809 230147 219843 230175
rect 219871 230147 235017 230175
rect 235045 230147 235079 230175
rect 235107 230147 235141 230175
rect 235169 230147 235203 230175
rect 235231 230147 250377 230175
rect 250405 230147 250439 230175
rect 250467 230147 250501 230175
rect 250529 230147 250563 230175
rect 250591 230147 265737 230175
rect 265765 230147 265799 230175
rect 265827 230147 265861 230175
rect 265889 230147 265923 230175
rect 265951 230147 281097 230175
rect 281125 230147 281159 230175
rect 281187 230147 281221 230175
rect 281249 230147 281283 230175
rect 281311 230147 296457 230175
rect 296485 230147 296519 230175
rect 296547 230147 296581 230175
rect 296609 230147 296643 230175
rect 296671 230147 298728 230175
rect 298756 230147 298790 230175
rect 298818 230147 298852 230175
rect 298880 230147 298914 230175
rect 298942 230147 298990 230175
rect -958 230113 298990 230147
rect -958 230085 -910 230113
rect -882 230085 -848 230113
rect -820 230085 -786 230113
rect -758 230085 -724 230113
rect -696 230085 4617 230113
rect 4645 230085 4679 230113
rect 4707 230085 4741 230113
rect 4769 230085 4803 230113
rect 4831 230085 29939 230113
rect 29967 230085 30001 230113
rect 30029 230085 45299 230113
rect 45327 230085 45361 230113
rect 45389 230085 60659 230113
rect 60687 230085 60721 230113
rect 60749 230085 76019 230113
rect 76047 230085 76081 230113
rect 76109 230085 96777 230113
rect 96805 230085 96839 230113
rect 96867 230085 96901 230113
rect 96929 230085 96963 230113
rect 96991 230085 109939 230113
rect 109967 230085 110001 230113
rect 110029 230085 125299 230113
rect 125327 230085 125361 230113
rect 125389 230085 140659 230113
rect 140687 230085 140721 230113
rect 140749 230085 156019 230113
rect 156047 230085 156081 230113
rect 156109 230085 173577 230113
rect 173605 230085 173639 230113
rect 173667 230085 173701 230113
rect 173729 230085 173763 230113
rect 173791 230085 188937 230113
rect 188965 230085 188999 230113
rect 189027 230085 189061 230113
rect 189089 230085 189123 230113
rect 189151 230085 204297 230113
rect 204325 230085 204359 230113
rect 204387 230085 204421 230113
rect 204449 230085 204483 230113
rect 204511 230085 219657 230113
rect 219685 230085 219719 230113
rect 219747 230085 219781 230113
rect 219809 230085 219843 230113
rect 219871 230085 235017 230113
rect 235045 230085 235079 230113
rect 235107 230085 235141 230113
rect 235169 230085 235203 230113
rect 235231 230085 250377 230113
rect 250405 230085 250439 230113
rect 250467 230085 250501 230113
rect 250529 230085 250563 230113
rect 250591 230085 265737 230113
rect 265765 230085 265799 230113
rect 265827 230085 265861 230113
rect 265889 230085 265923 230113
rect 265951 230085 281097 230113
rect 281125 230085 281159 230113
rect 281187 230085 281221 230113
rect 281249 230085 281283 230113
rect 281311 230085 296457 230113
rect 296485 230085 296519 230113
rect 296547 230085 296581 230113
rect 296609 230085 296643 230113
rect 296671 230085 298728 230113
rect 298756 230085 298790 230113
rect 298818 230085 298852 230113
rect 298880 230085 298914 230113
rect 298942 230085 298990 230113
rect -958 230051 298990 230085
rect -958 230023 -910 230051
rect -882 230023 -848 230051
rect -820 230023 -786 230051
rect -758 230023 -724 230051
rect -696 230023 4617 230051
rect 4645 230023 4679 230051
rect 4707 230023 4741 230051
rect 4769 230023 4803 230051
rect 4831 230023 29939 230051
rect 29967 230023 30001 230051
rect 30029 230023 45299 230051
rect 45327 230023 45361 230051
rect 45389 230023 60659 230051
rect 60687 230023 60721 230051
rect 60749 230023 76019 230051
rect 76047 230023 76081 230051
rect 76109 230023 96777 230051
rect 96805 230023 96839 230051
rect 96867 230023 96901 230051
rect 96929 230023 96963 230051
rect 96991 230023 109939 230051
rect 109967 230023 110001 230051
rect 110029 230023 125299 230051
rect 125327 230023 125361 230051
rect 125389 230023 140659 230051
rect 140687 230023 140721 230051
rect 140749 230023 156019 230051
rect 156047 230023 156081 230051
rect 156109 230023 173577 230051
rect 173605 230023 173639 230051
rect 173667 230023 173701 230051
rect 173729 230023 173763 230051
rect 173791 230023 188937 230051
rect 188965 230023 188999 230051
rect 189027 230023 189061 230051
rect 189089 230023 189123 230051
rect 189151 230023 204297 230051
rect 204325 230023 204359 230051
rect 204387 230023 204421 230051
rect 204449 230023 204483 230051
rect 204511 230023 219657 230051
rect 219685 230023 219719 230051
rect 219747 230023 219781 230051
rect 219809 230023 219843 230051
rect 219871 230023 235017 230051
rect 235045 230023 235079 230051
rect 235107 230023 235141 230051
rect 235169 230023 235203 230051
rect 235231 230023 250377 230051
rect 250405 230023 250439 230051
rect 250467 230023 250501 230051
rect 250529 230023 250563 230051
rect 250591 230023 265737 230051
rect 265765 230023 265799 230051
rect 265827 230023 265861 230051
rect 265889 230023 265923 230051
rect 265951 230023 281097 230051
rect 281125 230023 281159 230051
rect 281187 230023 281221 230051
rect 281249 230023 281283 230051
rect 281311 230023 296457 230051
rect 296485 230023 296519 230051
rect 296547 230023 296581 230051
rect 296609 230023 296643 230051
rect 296671 230023 298728 230051
rect 298756 230023 298790 230051
rect 298818 230023 298852 230051
rect 298880 230023 298914 230051
rect 298942 230023 298990 230051
rect -958 229989 298990 230023
rect -958 229961 -910 229989
rect -882 229961 -848 229989
rect -820 229961 -786 229989
rect -758 229961 -724 229989
rect -696 229961 4617 229989
rect 4645 229961 4679 229989
rect 4707 229961 4741 229989
rect 4769 229961 4803 229989
rect 4831 229961 29939 229989
rect 29967 229961 30001 229989
rect 30029 229961 45299 229989
rect 45327 229961 45361 229989
rect 45389 229961 60659 229989
rect 60687 229961 60721 229989
rect 60749 229961 76019 229989
rect 76047 229961 76081 229989
rect 76109 229961 96777 229989
rect 96805 229961 96839 229989
rect 96867 229961 96901 229989
rect 96929 229961 96963 229989
rect 96991 229961 109939 229989
rect 109967 229961 110001 229989
rect 110029 229961 125299 229989
rect 125327 229961 125361 229989
rect 125389 229961 140659 229989
rect 140687 229961 140721 229989
rect 140749 229961 156019 229989
rect 156047 229961 156081 229989
rect 156109 229961 173577 229989
rect 173605 229961 173639 229989
rect 173667 229961 173701 229989
rect 173729 229961 173763 229989
rect 173791 229961 188937 229989
rect 188965 229961 188999 229989
rect 189027 229961 189061 229989
rect 189089 229961 189123 229989
rect 189151 229961 204297 229989
rect 204325 229961 204359 229989
rect 204387 229961 204421 229989
rect 204449 229961 204483 229989
rect 204511 229961 219657 229989
rect 219685 229961 219719 229989
rect 219747 229961 219781 229989
rect 219809 229961 219843 229989
rect 219871 229961 235017 229989
rect 235045 229961 235079 229989
rect 235107 229961 235141 229989
rect 235169 229961 235203 229989
rect 235231 229961 250377 229989
rect 250405 229961 250439 229989
rect 250467 229961 250501 229989
rect 250529 229961 250563 229989
rect 250591 229961 265737 229989
rect 265765 229961 265799 229989
rect 265827 229961 265861 229989
rect 265889 229961 265923 229989
rect 265951 229961 281097 229989
rect 281125 229961 281159 229989
rect 281187 229961 281221 229989
rect 281249 229961 281283 229989
rect 281311 229961 296457 229989
rect 296485 229961 296519 229989
rect 296547 229961 296581 229989
rect 296609 229961 296643 229989
rect 296671 229961 298728 229989
rect 298756 229961 298790 229989
rect 298818 229961 298852 229989
rect 298880 229961 298914 229989
rect 298942 229961 298990 229989
rect -958 229913 298990 229961
rect -958 227175 298990 227223
rect -958 227147 -430 227175
rect -402 227147 -368 227175
rect -340 227147 -306 227175
rect -278 227147 -244 227175
rect -216 227147 2757 227175
rect 2785 227147 2819 227175
rect 2847 227147 2881 227175
rect 2909 227147 2943 227175
rect 2971 227147 18117 227175
rect 18145 227147 18179 227175
rect 18207 227147 18241 227175
rect 18269 227147 18303 227175
rect 18331 227147 22259 227175
rect 22287 227147 22321 227175
rect 22349 227147 37619 227175
rect 37647 227147 37681 227175
rect 37709 227147 52979 227175
rect 53007 227147 53041 227175
rect 53069 227147 68339 227175
rect 68367 227147 68401 227175
rect 68429 227147 83699 227175
rect 83727 227147 83761 227175
rect 83789 227147 94917 227175
rect 94945 227147 94979 227175
rect 95007 227147 95041 227175
rect 95069 227147 95103 227175
rect 95131 227147 102259 227175
rect 102287 227147 102321 227175
rect 102349 227147 117619 227175
rect 117647 227147 117681 227175
rect 117709 227147 132979 227175
rect 133007 227147 133041 227175
rect 133069 227147 148339 227175
rect 148367 227147 148401 227175
rect 148429 227147 163699 227175
rect 163727 227147 163761 227175
rect 163789 227147 171717 227175
rect 171745 227147 171779 227175
rect 171807 227147 171841 227175
rect 171869 227147 171903 227175
rect 171931 227147 187077 227175
rect 187105 227147 187139 227175
rect 187167 227147 187201 227175
rect 187229 227147 187263 227175
rect 187291 227147 202437 227175
rect 202465 227147 202499 227175
rect 202527 227147 202561 227175
rect 202589 227147 202623 227175
rect 202651 227147 217797 227175
rect 217825 227147 217859 227175
rect 217887 227147 217921 227175
rect 217949 227147 217983 227175
rect 218011 227147 233157 227175
rect 233185 227147 233219 227175
rect 233247 227147 233281 227175
rect 233309 227147 233343 227175
rect 233371 227147 248517 227175
rect 248545 227147 248579 227175
rect 248607 227147 248641 227175
rect 248669 227147 248703 227175
rect 248731 227147 263877 227175
rect 263905 227147 263939 227175
rect 263967 227147 264001 227175
rect 264029 227147 264063 227175
rect 264091 227147 279237 227175
rect 279265 227147 279299 227175
rect 279327 227147 279361 227175
rect 279389 227147 279423 227175
rect 279451 227147 294597 227175
rect 294625 227147 294659 227175
rect 294687 227147 294721 227175
rect 294749 227147 294783 227175
rect 294811 227147 298248 227175
rect 298276 227147 298310 227175
rect 298338 227147 298372 227175
rect 298400 227147 298434 227175
rect 298462 227147 298990 227175
rect -958 227113 298990 227147
rect -958 227085 -430 227113
rect -402 227085 -368 227113
rect -340 227085 -306 227113
rect -278 227085 -244 227113
rect -216 227085 2757 227113
rect 2785 227085 2819 227113
rect 2847 227085 2881 227113
rect 2909 227085 2943 227113
rect 2971 227085 18117 227113
rect 18145 227085 18179 227113
rect 18207 227085 18241 227113
rect 18269 227085 18303 227113
rect 18331 227085 22259 227113
rect 22287 227085 22321 227113
rect 22349 227085 37619 227113
rect 37647 227085 37681 227113
rect 37709 227085 52979 227113
rect 53007 227085 53041 227113
rect 53069 227085 68339 227113
rect 68367 227085 68401 227113
rect 68429 227085 83699 227113
rect 83727 227085 83761 227113
rect 83789 227085 94917 227113
rect 94945 227085 94979 227113
rect 95007 227085 95041 227113
rect 95069 227085 95103 227113
rect 95131 227085 102259 227113
rect 102287 227085 102321 227113
rect 102349 227085 117619 227113
rect 117647 227085 117681 227113
rect 117709 227085 132979 227113
rect 133007 227085 133041 227113
rect 133069 227085 148339 227113
rect 148367 227085 148401 227113
rect 148429 227085 163699 227113
rect 163727 227085 163761 227113
rect 163789 227085 171717 227113
rect 171745 227085 171779 227113
rect 171807 227085 171841 227113
rect 171869 227085 171903 227113
rect 171931 227085 187077 227113
rect 187105 227085 187139 227113
rect 187167 227085 187201 227113
rect 187229 227085 187263 227113
rect 187291 227085 202437 227113
rect 202465 227085 202499 227113
rect 202527 227085 202561 227113
rect 202589 227085 202623 227113
rect 202651 227085 217797 227113
rect 217825 227085 217859 227113
rect 217887 227085 217921 227113
rect 217949 227085 217983 227113
rect 218011 227085 233157 227113
rect 233185 227085 233219 227113
rect 233247 227085 233281 227113
rect 233309 227085 233343 227113
rect 233371 227085 248517 227113
rect 248545 227085 248579 227113
rect 248607 227085 248641 227113
rect 248669 227085 248703 227113
rect 248731 227085 263877 227113
rect 263905 227085 263939 227113
rect 263967 227085 264001 227113
rect 264029 227085 264063 227113
rect 264091 227085 279237 227113
rect 279265 227085 279299 227113
rect 279327 227085 279361 227113
rect 279389 227085 279423 227113
rect 279451 227085 294597 227113
rect 294625 227085 294659 227113
rect 294687 227085 294721 227113
rect 294749 227085 294783 227113
rect 294811 227085 298248 227113
rect 298276 227085 298310 227113
rect 298338 227085 298372 227113
rect 298400 227085 298434 227113
rect 298462 227085 298990 227113
rect -958 227051 298990 227085
rect -958 227023 -430 227051
rect -402 227023 -368 227051
rect -340 227023 -306 227051
rect -278 227023 -244 227051
rect -216 227023 2757 227051
rect 2785 227023 2819 227051
rect 2847 227023 2881 227051
rect 2909 227023 2943 227051
rect 2971 227023 18117 227051
rect 18145 227023 18179 227051
rect 18207 227023 18241 227051
rect 18269 227023 18303 227051
rect 18331 227023 22259 227051
rect 22287 227023 22321 227051
rect 22349 227023 37619 227051
rect 37647 227023 37681 227051
rect 37709 227023 52979 227051
rect 53007 227023 53041 227051
rect 53069 227023 68339 227051
rect 68367 227023 68401 227051
rect 68429 227023 83699 227051
rect 83727 227023 83761 227051
rect 83789 227023 94917 227051
rect 94945 227023 94979 227051
rect 95007 227023 95041 227051
rect 95069 227023 95103 227051
rect 95131 227023 102259 227051
rect 102287 227023 102321 227051
rect 102349 227023 117619 227051
rect 117647 227023 117681 227051
rect 117709 227023 132979 227051
rect 133007 227023 133041 227051
rect 133069 227023 148339 227051
rect 148367 227023 148401 227051
rect 148429 227023 163699 227051
rect 163727 227023 163761 227051
rect 163789 227023 171717 227051
rect 171745 227023 171779 227051
rect 171807 227023 171841 227051
rect 171869 227023 171903 227051
rect 171931 227023 187077 227051
rect 187105 227023 187139 227051
rect 187167 227023 187201 227051
rect 187229 227023 187263 227051
rect 187291 227023 202437 227051
rect 202465 227023 202499 227051
rect 202527 227023 202561 227051
rect 202589 227023 202623 227051
rect 202651 227023 217797 227051
rect 217825 227023 217859 227051
rect 217887 227023 217921 227051
rect 217949 227023 217983 227051
rect 218011 227023 233157 227051
rect 233185 227023 233219 227051
rect 233247 227023 233281 227051
rect 233309 227023 233343 227051
rect 233371 227023 248517 227051
rect 248545 227023 248579 227051
rect 248607 227023 248641 227051
rect 248669 227023 248703 227051
rect 248731 227023 263877 227051
rect 263905 227023 263939 227051
rect 263967 227023 264001 227051
rect 264029 227023 264063 227051
rect 264091 227023 279237 227051
rect 279265 227023 279299 227051
rect 279327 227023 279361 227051
rect 279389 227023 279423 227051
rect 279451 227023 294597 227051
rect 294625 227023 294659 227051
rect 294687 227023 294721 227051
rect 294749 227023 294783 227051
rect 294811 227023 298248 227051
rect 298276 227023 298310 227051
rect 298338 227023 298372 227051
rect 298400 227023 298434 227051
rect 298462 227023 298990 227051
rect -958 226989 298990 227023
rect -958 226961 -430 226989
rect -402 226961 -368 226989
rect -340 226961 -306 226989
rect -278 226961 -244 226989
rect -216 226961 2757 226989
rect 2785 226961 2819 226989
rect 2847 226961 2881 226989
rect 2909 226961 2943 226989
rect 2971 226961 18117 226989
rect 18145 226961 18179 226989
rect 18207 226961 18241 226989
rect 18269 226961 18303 226989
rect 18331 226961 22259 226989
rect 22287 226961 22321 226989
rect 22349 226961 37619 226989
rect 37647 226961 37681 226989
rect 37709 226961 52979 226989
rect 53007 226961 53041 226989
rect 53069 226961 68339 226989
rect 68367 226961 68401 226989
rect 68429 226961 83699 226989
rect 83727 226961 83761 226989
rect 83789 226961 94917 226989
rect 94945 226961 94979 226989
rect 95007 226961 95041 226989
rect 95069 226961 95103 226989
rect 95131 226961 102259 226989
rect 102287 226961 102321 226989
rect 102349 226961 117619 226989
rect 117647 226961 117681 226989
rect 117709 226961 132979 226989
rect 133007 226961 133041 226989
rect 133069 226961 148339 226989
rect 148367 226961 148401 226989
rect 148429 226961 163699 226989
rect 163727 226961 163761 226989
rect 163789 226961 171717 226989
rect 171745 226961 171779 226989
rect 171807 226961 171841 226989
rect 171869 226961 171903 226989
rect 171931 226961 187077 226989
rect 187105 226961 187139 226989
rect 187167 226961 187201 226989
rect 187229 226961 187263 226989
rect 187291 226961 202437 226989
rect 202465 226961 202499 226989
rect 202527 226961 202561 226989
rect 202589 226961 202623 226989
rect 202651 226961 217797 226989
rect 217825 226961 217859 226989
rect 217887 226961 217921 226989
rect 217949 226961 217983 226989
rect 218011 226961 233157 226989
rect 233185 226961 233219 226989
rect 233247 226961 233281 226989
rect 233309 226961 233343 226989
rect 233371 226961 248517 226989
rect 248545 226961 248579 226989
rect 248607 226961 248641 226989
rect 248669 226961 248703 226989
rect 248731 226961 263877 226989
rect 263905 226961 263939 226989
rect 263967 226961 264001 226989
rect 264029 226961 264063 226989
rect 264091 226961 279237 226989
rect 279265 226961 279299 226989
rect 279327 226961 279361 226989
rect 279389 226961 279423 226989
rect 279451 226961 294597 226989
rect 294625 226961 294659 226989
rect 294687 226961 294721 226989
rect 294749 226961 294783 226989
rect 294811 226961 298248 226989
rect 298276 226961 298310 226989
rect 298338 226961 298372 226989
rect 298400 226961 298434 226989
rect 298462 226961 298990 226989
rect -958 226913 298990 226961
rect -958 221175 298990 221223
rect -958 221147 -910 221175
rect -882 221147 -848 221175
rect -820 221147 -786 221175
rect -758 221147 -724 221175
rect -696 221147 4617 221175
rect 4645 221147 4679 221175
rect 4707 221147 4741 221175
rect 4769 221147 4803 221175
rect 4831 221147 29939 221175
rect 29967 221147 30001 221175
rect 30029 221147 45299 221175
rect 45327 221147 45361 221175
rect 45389 221147 60659 221175
rect 60687 221147 60721 221175
rect 60749 221147 76019 221175
rect 76047 221147 76081 221175
rect 76109 221147 96777 221175
rect 96805 221147 96839 221175
rect 96867 221147 96901 221175
rect 96929 221147 96963 221175
rect 96991 221147 109939 221175
rect 109967 221147 110001 221175
rect 110029 221147 125299 221175
rect 125327 221147 125361 221175
rect 125389 221147 140659 221175
rect 140687 221147 140721 221175
rect 140749 221147 156019 221175
rect 156047 221147 156081 221175
rect 156109 221147 173577 221175
rect 173605 221147 173639 221175
rect 173667 221147 173701 221175
rect 173729 221147 173763 221175
rect 173791 221147 188937 221175
rect 188965 221147 188999 221175
rect 189027 221147 189061 221175
rect 189089 221147 189123 221175
rect 189151 221147 204297 221175
rect 204325 221147 204359 221175
rect 204387 221147 204421 221175
rect 204449 221147 204483 221175
rect 204511 221147 219657 221175
rect 219685 221147 219719 221175
rect 219747 221147 219781 221175
rect 219809 221147 219843 221175
rect 219871 221147 235017 221175
rect 235045 221147 235079 221175
rect 235107 221147 235141 221175
rect 235169 221147 235203 221175
rect 235231 221147 250377 221175
rect 250405 221147 250439 221175
rect 250467 221147 250501 221175
rect 250529 221147 250563 221175
rect 250591 221147 265737 221175
rect 265765 221147 265799 221175
rect 265827 221147 265861 221175
rect 265889 221147 265923 221175
rect 265951 221147 281097 221175
rect 281125 221147 281159 221175
rect 281187 221147 281221 221175
rect 281249 221147 281283 221175
rect 281311 221147 296457 221175
rect 296485 221147 296519 221175
rect 296547 221147 296581 221175
rect 296609 221147 296643 221175
rect 296671 221147 298728 221175
rect 298756 221147 298790 221175
rect 298818 221147 298852 221175
rect 298880 221147 298914 221175
rect 298942 221147 298990 221175
rect -958 221113 298990 221147
rect -958 221085 -910 221113
rect -882 221085 -848 221113
rect -820 221085 -786 221113
rect -758 221085 -724 221113
rect -696 221085 4617 221113
rect 4645 221085 4679 221113
rect 4707 221085 4741 221113
rect 4769 221085 4803 221113
rect 4831 221085 29939 221113
rect 29967 221085 30001 221113
rect 30029 221085 45299 221113
rect 45327 221085 45361 221113
rect 45389 221085 60659 221113
rect 60687 221085 60721 221113
rect 60749 221085 76019 221113
rect 76047 221085 76081 221113
rect 76109 221085 96777 221113
rect 96805 221085 96839 221113
rect 96867 221085 96901 221113
rect 96929 221085 96963 221113
rect 96991 221085 109939 221113
rect 109967 221085 110001 221113
rect 110029 221085 125299 221113
rect 125327 221085 125361 221113
rect 125389 221085 140659 221113
rect 140687 221085 140721 221113
rect 140749 221085 156019 221113
rect 156047 221085 156081 221113
rect 156109 221085 173577 221113
rect 173605 221085 173639 221113
rect 173667 221085 173701 221113
rect 173729 221085 173763 221113
rect 173791 221085 188937 221113
rect 188965 221085 188999 221113
rect 189027 221085 189061 221113
rect 189089 221085 189123 221113
rect 189151 221085 204297 221113
rect 204325 221085 204359 221113
rect 204387 221085 204421 221113
rect 204449 221085 204483 221113
rect 204511 221085 219657 221113
rect 219685 221085 219719 221113
rect 219747 221085 219781 221113
rect 219809 221085 219843 221113
rect 219871 221085 235017 221113
rect 235045 221085 235079 221113
rect 235107 221085 235141 221113
rect 235169 221085 235203 221113
rect 235231 221085 250377 221113
rect 250405 221085 250439 221113
rect 250467 221085 250501 221113
rect 250529 221085 250563 221113
rect 250591 221085 265737 221113
rect 265765 221085 265799 221113
rect 265827 221085 265861 221113
rect 265889 221085 265923 221113
rect 265951 221085 281097 221113
rect 281125 221085 281159 221113
rect 281187 221085 281221 221113
rect 281249 221085 281283 221113
rect 281311 221085 296457 221113
rect 296485 221085 296519 221113
rect 296547 221085 296581 221113
rect 296609 221085 296643 221113
rect 296671 221085 298728 221113
rect 298756 221085 298790 221113
rect 298818 221085 298852 221113
rect 298880 221085 298914 221113
rect 298942 221085 298990 221113
rect -958 221051 298990 221085
rect -958 221023 -910 221051
rect -882 221023 -848 221051
rect -820 221023 -786 221051
rect -758 221023 -724 221051
rect -696 221023 4617 221051
rect 4645 221023 4679 221051
rect 4707 221023 4741 221051
rect 4769 221023 4803 221051
rect 4831 221023 29939 221051
rect 29967 221023 30001 221051
rect 30029 221023 45299 221051
rect 45327 221023 45361 221051
rect 45389 221023 60659 221051
rect 60687 221023 60721 221051
rect 60749 221023 76019 221051
rect 76047 221023 76081 221051
rect 76109 221023 96777 221051
rect 96805 221023 96839 221051
rect 96867 221023 96901 221051
rect 96929 221023 96963 221051
rect 96991 221023 109939 221051
rect 109967 221023 110001 221051
rect 110029 221023 125299 221051
rect 125327 221023 125361 221051
rect 125389 221023 140659 221051
rect 140687 221023 140721 221051
rect 140749 221023 156019 221051
rect 156047 221023 156081 221051
rect 156109 221023 173577 221051
rect 173605 221023 173639 221051
rect 173667 221023 173701 221051
rect 173729 221023 173763 221051
rect 173791 221023 188937 221051
rect 188965 221023 188999 221051
rect 189027 221023 189061 221051
rect 189089 221023 189123 221051
rect 189151 221023 204297 221051
rect 204325 221023 204359 221051
rect 204387 221023 204421 221051
rect 204449 221023 204483 221051
rect 204511 221023 219657 221051
rect 219685 221023 219719 221051
rect 219747 221023 219781 221051
rect 219809 221023 219843 221051
rect 219871 221023 235017 221051
rect 235045 221023 235079 221051
rect 235107 221023 235141 221051
rect 235169 221023 235203 221051
rect 235231 221023 250377 221051
rect 250405 221023 250439 221051
rect 250467 221023 250501 221051
rect 250529 221023 250563 221051
rect 250591 221023 265737 221051
rect 265765 221023 265799 221051
rect 265827 221023 265861 221051
rect 265889 221023 265923 221051
rect 265951 221023 281097 221051
rect 281125 221023 281159 221051
rect 281187 221023 281221 221051
rect 281249 221023 281283 221051
rect 281311 221023 296457 221051
rect 296485 221023 296519 221051
rect 296547 221023 296581 221051
rect 296609 221023 296643 221051
rect 296671 221023 298728 221051
rect 298756 221023 298790 221051
rect 298818 221023 298852 221051
rect 298880 221023 298914 221051
rect 298942 221023 298990 221051
rect -958 220989 298990 221023
rect -958 220961 -910 220989
rect -882 220961 -848 220989
rect -820 220961 -786 220989
rect -758 220961 -724 220989
rect -696 220961 4617 220989
rect 4645 220961 4679 220989
rect 4707 220961 4741 220989
rect 4769 220961 4803 220989
rect 4831 220961 29939 220989
rect 29967 220961 30001 220989
rect 30029 220961 45299 220989
rect 45327 220961 45361 220989
rect 45389 220961 60659 220989
rect 60687 220961 60721 220989
rect 60749 220961 76019 220989
rect 76047 220961 76081 220989
rect 76109 220961 96777 220989
rect 96805 220961 96839 220989
rect 96867 220961 96901 220989
rect 96929 220961 96963 220989
rect 96991 220961 109939 220989
rect 109967 220961 110001 220989
rect 110029 220961 125299 220989
rect 125327 220961 125361 220989
rect 125389 220961 140659 220989
rect 140687 220961 140721 220989
rect 140749 220961 156019 220989
rect 156047 220961 156081 220989
rect 156109 220961 173577 220989
rect 173605 220961 173639 220989
rect 173667 220961 173701 220989
rect 173729 220961 173763 220989
rect 173791 220961 188937 220989
rect 188965 220961 188999 220989
rect 189027 220961 189061 220989
rect 189089 220961 189123 220989
rect 189151 220961 204297 220989
rect 204325 220961 204359 220989
rect 204387 220961 204421 220989
rect 204449 220961 204483 220989
rect 204511 220961 219657 220989
rect 219685 220961 219719 220989
rect 219747 220961 219781 220989
rect 219809 220961 219843 220989
rect 219871 220961 235017 220989
rect 235045 220961 235079 220989
rect 235107 220961 235141 220989
rect 235169 220961 235203 220989
rect 235231 220961 250377 220989
rect 250405 220961 250439 220989
rect 250467 220961 250501 220989
rect 250529 220961 250563 220989
rect 250591 220961 265737 220989
rect 265765 220961 265799 220989
rect 265827 220961 265861 220989
rect 265889 220961 265923 220989
rect 265951 220961 281097 220989
rect 281125 220961 281159 220989
rect 281187 220961 281221 220989
rect 281249 220961 281283 220989
rect 281311 220961 296457 220989
rect 296485 220961 296519 220989
rect 296547 220961 296581 220989
rect 296609 220961 296643 220989
rect 296671 220961 298728 220989
rect 298756 220961 298790 220989
rect 298818 220961 298852 220989
rect 298880 220961 298914 220989
rect 298942 220961 298990 220989
rect -958 220913 298990 220961
rect -958 218175 298990 218223
rect -958 218147 -430 218175
rect -402 218147 -368 218175
rect -340 218147 -306 218175
rect -278 218147 -244 218175
rect -216 218147 2757 218175
rect 2785 218147 2819 218175
rect 2847 218147 2881 218175
rect 2909 218147 2943 218175
rect 2971 218147 18117 218175
rect 18145 218147 18179 218175
rect 18207 218147 18241 218175
rect 18269 218147 18303 218175
rect 18331 218147 22259 218175
rect 22287 218147 22321 218175
rect 22349 218147 37619 218175
rect 37647 218147 37681 218175
rect 37709 218147 52979 218175
rect 53007 218147 53041 218175
rect 53069 218147 68339 218175
rect 68367 218147 68401 218175
rect 68429 218147 83699 218175
rect 83727 218147 83761 218175
rect 83789 218147 94917 218175
rect 94945 218147 94979 218175
rect 95007 218147 95041 218175
rect 95069 218147 95103 218175
rect 95131 218147 102259 218175
rect 102287 218147 102321 218175
rect 102349 218147 117619 218175
rect 117647 218147 117681 218175
rect 117709 218147 132979 218175
rect 133007 218147 133041 218175
rect 133069 218147 148339 218175
rect 148367 218147 148401 218175
rect 148429 218147 163699 218175
rect 163727 218147 163761 218175
rect 163789 218147 171717 218175
rect 171745 218147 171779 218175
rect 171807 218147 171841 218175
rect 171869 218147 171903 218175
rect 171931 218147 187077 218175
rect 187105 218147 187139 218175
rect 187167 218147 187201 218175
rect 187229 218147 187263 218175
rect 187291 218147 202437 218175
rect 202465 218147 202499 218175
rect 202527 218147 202561 218175
rect 202589 218147 202623 218175
rect 202651 218147 217797 218175
rect 217825 218147 217859 218175
rect 217887 218147 217921 218175
rect 217949 218147 217983 218175
rect 218011 218147 233157 218175
rect 233185 218147 233219 218175
rect 233247 218147 233281 218175
rect 233309 218147 233343 218175
rect 233371 218147 248517 218175
rect 248545 218147 248579 218175
rect 248607 218147 248641 218175
rect 248669 218147 248703 218175
rect 248731 218147 263877 218175
rect 263905 218147 263939 218175
rect 263967 218147 264001 218175
rect 264029 218147 264063 218175
rect 264091 218147 279237 218175
rect 279265 218147 279299 218175
rect 279327 218147 279361 218175
rect 279389 218147 279423 218175
rect 279451 218147 294597 218175
rect 294625 218147 294659 218175
rect 294687 218147 294721 218175
rect 294749 218147 294783 218175
rect 294811 218147 298248 218175
rect 298276 218147 298310 218175
rect 298338 218147 298372 218175
rect 298400 218147 298434 218175
rect 298462 218147 298990 218175
rect -958 218113 298990 218147
rect -958 218085 -430 218113
rect -402 218085 -368 218113
rect -340 218085 -306 218113
rect -278 218085 -244 218113
rect -216 218085 2757 218113
rect 2785 218085 2819 218113
rect 2847 218085 2881 218113
rect 2909 218085 2943 218113
rect 2971 218085 18117 218113
rect 18145 218085 18179 218113
rect 18207 218085 18241 218113
rect 18269 218085 18303 218113
rect 18331 218085 22259 218113
rect 22287 218085 22321 218113
rect 22349 218085 37619 218113
rect 37647 218085 37681 218113
rect 37709 218085 52979 218113
rect 53007 218085 53041 218113
rect 53069 218085 68339 218113
rect 68367 218085 68401 218113
rect 68429 218085 83699 218113
rect 83727 218085 83761 218113
rect 83789 218085 94917 218113
rect 94945 218085 94979 218113
rect 95007 218085 95041 218113
rect 95069 218085 95103 218113
rect 95131 218085 102259 218113
rect 102287 218085 102321 218113
rect 102349 218085 117619 218113
rect 117647 218085 117681 218113
rect 117709 218085 132979 218113
rect 133007 218085 133041 218113
rect 133069 218085 148339 218113
rect 148367 218085 148401 218113
rect 148429 218085 163699 218113
rect 163727 218085 163761 218113
rect 163789 218085 171717 218113
rect 171745 218085 171779 218113
rect 171807 218085 171841 218113
rect 171869 218085 171903 218113
rect 171931 218085 187077 218113
rect 187105 218085 187139 218113
rect 187167 218085 187201 218113
rect 187229 218085 187263 218113
rect 187291 218085 202437 218113
rect 202465 218085 202499 218113
rect 202527 218085 202561 218113
rect 202589 218085 202623 218113
rect 202651 218085 217797 218113
rect 217825 218085 217859 218113
rect 217887 218085 217921 218113
rect 217949 218085 217983 218113
rect 218011 218085 233157 218113
rect 233185 218085 233219 218113
rect 233247 218085 233281 218113
rect 233309 218085 233343 218113
rect 233371 218085 248517 218113
rect 248545 218085 248579 218113
rect 248607 218085 248641 218113
rect 248669 218085 248703 218113
rect 248731 218085 263877 218113
rect 263905 218085 263939 218113
rect 263967 218085 264001 218113
rect 264029 218085 264063 218113
rect 264091 218085 279237 218113
rect 279265 218085 279299 218113
rect 279327 218085 279361 218113
rect 279389 218085 279423 218113
rect 279451 218085 294597 218113
rect 294625 218085 294659 218113
rect 294687 218085 294721 218113
rect 294749 218085 294783 218113
rect 294811 218085 298248 218113
rect 298276 218085 298310 218113
rect 298338 218085 298372 218113
rect 298400 218085 298434 218113
rect 298462 218085 298990 218113
rect -958 218051 298990 218085
rect -958 218023 -430 218051
rect -402 218023 -368 218051
rect -340 218023 -306 218051
rect -278 218023 -244 218051
rect -216 218023 2757 218051
rect 2785 218023 2819 218051
rect 2847 218023 2881 218051
rect 2909 218023 2943 218051
rect 2971 218023 18117 218051
rect 18145 218023 18179 218051
rect 18207 218023 18241 218051
rect 18269 218023 18303 218051
rect 18331 218023 22259 218051
rect 22287 218023 22321 218051
rect 22349 218023 37619 218051
rect 37647 218023 37681 218051
rect 37709 218023 52979 218051
rect 53007 218023 53041 218051
rect 53069 218023 68339 218051
rect 68367 218023 68401 218051
rect 68429 218023 83699 218051
rect 83727 218023 83761 218051
rect 83789 218023 94917 218051
rect 94945 218023 94979 218051
rect 95007 218023 95041 218051
rect 95069 218023 95103 218051
rect 95131 218023 102259 218051
rect 102287 218023 102321 218051
rect 102349 218023 117619 218051
rect 117647 218023 117681 218051
rect 117709 218023 132979 218051
rect 133007 218023 133041 218051
rect 133069 218023 148339 218051
rect 148367 218023 148401 218051
rect 148429 218023 163699 218051
rect 163727 218023 163761 218051
rect 163789 218023 171717 218051
rect 171745 218023 171779 218051
rect 171807 218023 171841 218051
rect 171869 218023 171903 218051
rect 171931 218023 187077 218051
rect 187105 218023 187139 218051
rect 187167 218023 187201 218051
rect 187229 218023 187263 218051
rect 187291 218023 202437 218051
rect 202465 218023 202499 218051
rect 202527 218023 202561 218051
rect 202589 218023 202623 218051
rect 202651 218023 217797 218051
rect 217825 218023 217859 218051
rect 217887 218023 217921 218051
rect 217949 218023 217983 218051
rect 218011 218023 233157 218051
rect 233185 218023 233219 218051
rect 233247 218023 233281 218051
rect 233309 218023 233343 218051
rect 233371 218023 248517 218051
rect 248545 218023 248579 218051
rect 248607 218023 248641 218051
rect 248669 218023 248703 218051
rect 248731 218023 263877 218051
rect 263905 218023 263939 218051
rect 263967 218023 264001 218051
rect 264029 218023 264063 218051
rect 264091 218023 279237 218051
rect 279265 218023 279299 218051
rect 279327 218023 279361 218051
rect 279389 218023 279423 218051
rect 279451 218023 294597 218051
rect 294625 218023 294659 218051
rect 294687 218023 294721 218051
rect 294749 218023 294783 218051
rect 294811 218023 298248 218051
rect 298276 218023 298310 218051
rect 298338 218023 298372 218051
rect 298400 218023 298434 218051
rect 298462 218023 298990 218051
rect -958 217989 298990 218023
rect -958 217961 -430 217989
rect -402 217961 -368 217989
rect -340 217961 -306 217989
rect -278 217961 -244 217989
rect -216 217961 2757 217989
rect 2785 217961 2819 217989
rect 2847 217961 2881 217989
rect 2909 217961 2943 217989
rect 2971 217961 18117 217989
rect 18145 217961 18179 217989
rect 18207 217961 18241 217989
rect 18269 217961 18303 217989
rect 18331 217961 22259 217989
rect 22287 217961 22321 217989
rect 22349 217961 37619 217989
rect 37647 217961 37681 217989
rect 37709 217961 52979 217989
rect 53007 217961 53041 217989
rect 53069 217961 68339 217989
rect 68367 217961 68401 217989
rect 68429 217961 83699 217989
rect 83727 217961 83761 217989
rect 83789 217961 94917 217989
rect 94945 217961 94979 217989
rect 95007 217961 95041 217989
rect 95069 217961 95103 217989
rect 95131 217961 102259 217989
rect 102287 217961 102321 217989
rect 102349 217961 117619 217989
rect 117647 217961 117681 217989
rect 117709 217961 132979 217989
rect 133007 217961 133041 217989
rect 133069 217961 148339 217989
rect 148367 217961 148401 217989
rect 148429 217961 163699 217989
rect 163727 217961 163761 217989
rect 163789 217961 171717 217989
rect 171745 217961 171779 217989
rect 171807 217961 171841 217989
rect 171869 217961 171903 217989
rect 171931 217961 187077 217989
rect 187105 217961 187139 217989
rect 187167 217961 187201 217989
rect 187229 217961 187263 217989
rect 187291 217961 202437 217989
rect 202465 217961 202499 217989
rect 202527 217961 202561 217989
rect 202589 217961 202623 217989
rect 202651 217961 217797 217989
rect 217825 217961 217859 217989
rect 217887 217961 217921 217989
rect 217949 217961 217983 217989
rect 218011 217961 233157 217989
rect 233185 217961 233219 217989
rect 233247 217961 233281 217989
rect 233309 217961 233343 217989
rect 233371 217961 248517 217989
rect 248545 217961 248579 217989
rect 248607 217961 248641 217989
rect 248669 217961 248703 217989
rect 248731 217961 263877 217989
rect 263905 217961 263939 217989
rect 263967 217961 264001 217989
rect 264029 217961 264063 217989
rect 264091 217961 279237 217989
rect 279265 217961 279299 217989
rect 279327 217961 279361 217989
rect 279389 217961 279423 217989
rect 279451 217961 294597 217989
rect 294625 217961 294659 217989
rect 294687 217961 294721 217989
rect 294749 217961 294783 217989
rect 294811 217961 298248 217989
rect 298276 217961 298310 217989
rect 298338 217961 298372 217989
rect 298400 217961 298434 217989
rect 298462 217961 298990 217989
rect -958 217913 298990 217961
rect -958 212175 298990 212223
rect -958 212147 -910 212175
rect -882 212147 -848 212175
rect -820 212147 -786 212175
rect -758 212147 -724 212175
rect -696 212147 4617 212175
rect 4645 212147 4679 212175
rect 4707 212147 4741 212175
rect 4769 212147 4803 212175
rect 4831 212147 29939 212175
rect 29967 212147 30001 212175
rect 30029 212147 45299 212175
rect 45327 212147 45361 212175
rect 45389 212147 60659 212175
rect 60687 212147 60721 212175
rect 60749 212147 76019 212175
rect 76047 212147 76081 212175
rect 76109 212147 96777 212175
rect 96805 212147 96839 212175
rect 96867 212147 96901 212175
rect 96929 212147 96963 212175
rect 96991 212147 109939 212175
rect 109967 212147 110001 212175
rect 110029 212147 125299 212175
rect 125327 212147 125361 212175
rect 125389 212147 140659 212175
rect 140687 212147 140721 212175
rect 140749 212147 156019 212175
rect 156047 212147 156081 212175
rect 156109 212147 173577 212175
rect 173605 212147 173639 212175
rect 173667 212147 173701 212175
rect 173729 212147 173763 212175
rect 173791 212147 188937 212175
rect 188965 212147 188999 212175
rect 189027 212147 189061 212175
rect 189089 212147 189123 212175
rect 189151 212147 204297 212175
rect 204325 212147 204359 212175
rect 204387 212147 204421 212175
rect 204449 212147 204483 212175
rect 204511 212147 219657 212175
rect 219685 212147 219719 212175
rect 219747 212147 219781 212175
rect 219809 212147 219843 212175
rect 219871 212147 235017 212175
rect 235045 212147 235079 212175
rect 235107 212147 235141 212175
rect 235169 212147 235203 212175
rect 235231 212147 250377 212175
rect 250405 212147 250439 212175
rect 250467 212147 250501 212175
rect 250529 212147 250563 212175
rect 250591 212147 265737 212175
rect 265765 212147 265799 212175
rect 265827 212147 265861 212175
rect 265889 212147 265923 212175
rect 265951 212147 281097 212175
rect 281125 212147 281159 212175
rect 281187 212147 281221 212175
rect 281249 212147 281283 212175
rect 281311 212147 296457 212175
rect 296485 212147 296519 212175
rect 296547 212147 296581 212175
rect 296609 212147 296643 212175
rect 296671 212147 298728 212175
rect 298756 212147 298790 212175
rect 298818 212147 298852 212175
rect 298880 212147 298914 212175
rect 298942 212147 298990 212175
rect -958 212113 298990 212147
rect -958 212085 -910 212113
rect -882 212085 -848 212113
rect -820 212085 -786 212113
rect -758 212085 -724 212113
rect -696 212085 4617 212113
rect 4645 212085 4679 212113
rect 4707 212085 4741 212113
rect 4769 212085 4803 212113
rect 4831 212085 29939 212113
rect 29967 212085 30001 212113
rect 30029 212085 45299 212113
rect 45327 212085 45361 212113
rect 45389 212085 60659 212113
rect 60687 212085 60721 212113
rect 60749 212085 76019 212113
rect 76047 212085 76081 212113
rect 76109 212085 96777 212113
rect 96805 212085 96839 212113
rect 96867 212085 96901 212113
rect 96929 212085 96963 212113
rect 96991 212085 109939 212113
rect 109967 212085 110001 212113
rect 110029 212085 125299 212113
rect 125327 212085 125361 212113
rect 125389 212085 140659 212113
rect 140687 212085 140721 212113
rect 140749 212085 156019 212113
rect 156047 212085 156081 212113
rect 156109 212085 173577 212113
rect 173605 212085 173639 212113
rect 173667 212085 173701 212113
rect 173729 212085 173763 212113
rect 173791 212085 188937 212113
rect 188965 212085 188999 212113
rect 189027 212085 189061 212113
rect 189089 212085 189123 212113
rect 189151 212085 204297 212113
rect 204325 212085 204359 212113
rect 204387 212085 204421 212113
rect 204449 212085 204483 212113
rect 204511 212085 219657 212113
rect 219685 212085 219719 212113
rect 219747 212085 219781 212113
rect 219809 212085 219843 212113
rect 219871 212085 235017 212113
rect 235045 212085 235079 212113
rect 235107 212085 235141 212113
rect 235169 212085 235203 212113
rect 235231 212085 250377 212113
rect 250405 212085 250439 212113
rect 250467 212085 250501 212113
rect 250529 212085 250563 212113
rect 250591 212085 265737 212113
rect 265765 212085 265799 212113
rect 265827 212085 265861 212113
rect 265889 212085 265923 212113
rect 265951 212085 281097 212113
rect 281125 212085 281159 212113
rect 281187 212085 281221 212113
rect 281249 212085 281283 212113
rect 281311 212085 296457 212113
rect 296485 212085 296519 212113
rect 296547 212085 296581 212113
rect 296609 212085 296643 212113
rect 296671 212085 298728 212113
rect 298756 212085 298790 212113
rect 298818 212085 298852 212113
rect 298880 212085 298914 212113
rect 298942 212085 298990 212113
rect -958 212051 298990 212085
rect -958 212023 -910 212051
rect -882 212023 -848 212051
rect -820 212023 -786 212051
rect -758 212023 -724 212051
rect -696 212023 4617 212051
rect 4645 212023 4679 212051
rect 4707 212023 4741 212051
rect 4769 212023 4803 212051
rect 4831 212023 29939 212051
rect 29967 212023 30001 212051
rect 30029 212023 45299 212051
rect 45327 212023 45361 212051
rect 45389 212023 60659 212051
rect 60687 212023 60721 212051
rect 60749 212023 76019 212051
rect 76047 212023 76081 212051
rect 76109 212023 96777 212051
rect 96805 212023 96839 212051
rect 96867 212023 96901 212051
rect 96929 212023 96963 212051
rect 96991 212023 109939 212051
rect 109967 212023 110001 212051
rect 110029 212023 125299 212051
rect 125327 212023 125361 212051
rect 125389 212023 140659 212051
rect 140687 212023 140721 212051
rect 140749 212023 156019 212051
rect 156047 212023 156081 212051
rect 156109 212023 173577 212051
rect 173605 212023 173639 212051
rect 173667 212023 173701 212051
rect 173729 212023 173763 212051
rect 173791 212023 188937 212051
rect 188965 212023 188999 212051
rect 189027 212023 189061 212051
rect 189089 212023 189123 212051
rect 189151 212023 204297 212051
rect 204325 212023 204359 212051
rect 204387 212023 204421 212051
rect 204449 212023 204483 212051
rect 204511 212023 219657 212051
rect 219685 212023 219719 212051
rect 219747 212023 219781 212051
rect 219809 212023 219843 212051
rect 219871 212023 235017 212051
rect 235045 212023 235079 212051
rect 235107 212023 235141 212051
rect 235169 212023 235203 212051
rect 235231 212023 250377 212051
rect 250405 212023 250439 212051
rect 250467 212023 250501 212051
rect 250529 212023 250563 212051
rect 250591 212023 265737 212051
rect 265765 212023 265799 212051
rect 265827 212023 265861 212051
rect 265889 212023 265923 212051
rect 265951 212023 281097 212051
rect 281125 212023 281159 212051
rect 281187 212023 281221 212051
rect 281249 212023 281283 212051
rect 281311 212023 296457 212051
rect 296485 212023 296519 212051
rect 296547 212023 296581 212051
rect 296609 212023 296643 212051
rect 296671 212023 298728 212051
rect 298756 212023 298790 212051
rect 298818 212023 298852 212051
rect 298880 212023 298914 212051
rect 298942 212023 298990 212051
rect -958 211989 298990 212023
rect -958 211961 -910 211989
rect -882 211961 -848 211989
rect -820 211961 -786 211989
rect -758 211961 -724 211989
rect -696 211961 4617 211989
rect 4645 211961 4679 211989
rect 4707 211961 4741 211989
rect 4769 211961 4803 211989
rect 4831 211961 29939 211989
rect 29967 211961 30001 211989
rect 30029 211961 45299 211989
rect 45327 211961 45361 211989
rect 45389 211961 60659 211989
rect 60687 211961 60721 211989
rect 60749 211961 76019 211989
rect 76047 211961 76081 211989
rect 76109 211961 96777 211989
rect 96805 211961 96839 211989
rect 96867 211961 96901 211989
rect 96929 211961 96963 211989
rect 96991 211961 109939 211989
rect 109967 211961 110001 211989
rect 110029 211961 125299 211989
rect 125327 211961 125361 211989
rect 125389 211961 140659 211989
rect 140687 211961 140721 211989
rect 140749 211961 156019 211989
rect 156047 211961 156081 211989
rect 156109 211961 173577 211989
rect 173605 211961 173639 211989
rect 173667 211961 173701 211989
rect 173729 211961 173763 211989
rect 173791 211961 188937 211989
rect 188965 211961 188999 211989
rect 189027 211961 189061 211989
rect 189089 211961 189123 211989
rect 189151 211961 204297 211989
rect 204325 211961 204359 211989
rect 204387 211961 204421 211989
rect 204449 211961 204483 211989
rect 204511 211961 219657 211989
rect 219685 211961 219719 211989
rect 219747 211961 219781 211989
rect 219809 211961 219843 211989
rect 219871 211961 235017 211989
rect 235045 211961 235079 211989
rect 235107 211961 235141 211989
rect 235169 211961 235203 211989
rect 235231 211961 250377 211989
rect 250405 211961 250439 211989
rect 250467 211961 250501 211989
rect 250529 211961 250563 211989
rect 250591 211961 265737 211989
rect 265765 211961 265799 211989
rect 265827 211961 265861 211989
rect 265889 211961 265923 211989
rect 265951 211961 281097 211989
rect 281125 211961 281159 211989
rect 281187 211961 281221 211989
rect 281249 211961 281283 211989
rect 281311 211961 296457 211989
rect 296485 211961 296519 211989
rect 296547 211961 296581 211989
rect 296609 211961 296643 211989
rect 296671 211961 298728 211989
rect 298756 211961 298790 211989
rect 298818 211961 298852 211989
rect 298880 211961 298914 211989
rect 298942 211961 298990 211989
rect -958 211913 298990 211961
rect -958 209175 298990 209223
rect -958 209147 -430 209175
rect -402 209147 -368 209175
rect -340 209147 -306 209175
rect -278 209147 -244 209175
rect -216 209147 2757 209175
rect 2785 209147 2819 209175
rect 2847 209147 2881 209175
rect 2909 209147 2943 209175
rect 2971 209147 18117 209175
rect 18145 209147 18179 209175
rect 18207 209147 18241 209175
rect 18269 209147 18303 209175
rect 18331 209147 22259 209175
rect 22287 209147 22321 209175
rect 22349 209147 37619 209175
rect 37647 209147 37681 209175
rect 37709 209147 52979 209175
rect 53007 209147 53041 209175
rect 53069 209147 68339 209175
rect 68367 209147 68401 209175
rect 68429 209147 83699 209175
rect 83727 209147 83761 209175
rect 83789 209147 94917 209175
rect 94945 209147 94979 209175
rect 95007 209147 95041 209175
rect 95069 209147 95103 209175
rect 95131 209147 102259 209175
rect 102287 209147 102321 209175
rect 102349 209147 117619 209175
rect 117647 209147 117681 209175
rect 117709 209147 132979 209175
rect 133007 209147 133041 209175
rect 133069 209147 148339 209175
rect 148367 209147 148401 209175
rect 148429 209147 163699 209175
rect 163727 209147 163761 209175
rect 163789 209147 171717 209175
rect 171745 209147 171779 209175
rect 171807 209147 171841 209175
rect 171869 209147 171903 209175
rect 171931 209147 187077 209175
rect 187105 209147 187139 209175
rect 187167 209147 187201 209175
rect 187229 209147 187263 209175
rect 187291 209147 202437 209175
rect 202465 209147 202499 209175
rect 202527 209147 202561 209175
rect 202589 209147 202623 209175
rect 202651 209147 217797 209175
rect 217825 209147 217859 209175
rect 217887 209147 217921 209175
rect 217949 209147 217983 209175
rect 218011 209147 233157 209175
rect 233185 209147 233219 209175
rect 233247 209147 233281 209175
rect 233309 209147 233343 209175
rect 233371 209147 248517 209175
rect 248545 209147 248579 209175
rect 248607 209147 248641 209175
rect 248669 209147 248703 209175
rect 248731 209147 263877 209175
rect 263905 209147 263939 209175
rect 263967 209147 264001 209175
rect 264029 209147 264063 209175
rect 264091 209147 279237 209175
rect 279265 209147 279299 209175
rect 279327 209147 279361 209175
rect 279389 209147 279423 209175
rect 279451 209147 294597 209175
rect 294625 209147 294659 209175
rect 294687 209147 294721 209175
rect 294749 209147 294783 209175
rect 294811 209147 298248 209175
rect 298276 209147 298310 209175
rect 298338 209147 298372 209175
rect 298400 209147 298434 209175
rect 298462 209147 298990 209175
rect -958 209113 298990 209147
rect -958 209085 -430 209113
rect -402 209085 -368 209113
rect -340 209085 -306 209113
rect -278 209085 -244 209113
rect -216 209085 2757 209113
rect 2785 209085 2819 209113
rect 2847 209085 2881 209113
rect 2909 209085 2943 209113
rect 2971 209085 18117 209113
rect 18145 209085 18179 209113
rect 18207 209085 18241 209113
rect 18269 209085 18303 209113
rect 18331 209085 22259 209113
rect 22287 209085 22321 209113
rect 22349 209085 37619 209113
rect 37647 209085 37681 209113
rect 37709 209085 52979 209113
rect 53007 209085 53041 209113
rect 53069 209085 68339 209113
rect 68367 209085 68401 209113
rect 68429 209085 83699 209113
rect 83727 209085 83761 209113
rect 83789 209085 94917 209113
rect 94945 209085 94979 209113
rect 95007 209085 95041 209113
rect 95069 209085 95103 209113
rect 95131 209085 102259 209113
rect 102287 209085 102321 209113
rect 102349 209085 117619 209113
rect 117647 209085 117681 209113
rect 117709 209085 132979 209113
rect 133007 209085 133041 209113
rect 133069 209085 148339 209113
rect 148367 209085 148401 209113
rect 148429 209085 163699 209113
rect 163727 209085 163761 209113
rect 163789 209085 171717 209113
rect 171745 209085 171779 209113
rect 171807 209085 171841 209113
rect 171869 209085 171903 209113
rect 171931 209085 187077 209113
rect 187105 209085 187139 209113
rect 187167 209085 187201 209113
rect 187229 209085 187263 209113
rect 187291 209085 202437 209113
rect 202465 209085 202499 209113
rect 202527 209085 202561 209113
rect 202589 209085 202623 209113
rect 202651 209085 217797 209113
rect 217825 209085 217859 209113
rect 217887 209085 217921 209113
rect 217949 209085 217983 209113
rect 218011 209085 233157 209113
rect 233185 209085 233219 209113
rect 233247 209085 233281 209113
rect 233309 209085 233343 209113
rect 233371 209085 248517 209113
rect 248545 209085 248579 209113
rect 248607 209085 248641 209113
rect 248669 209085 248703 209113
rect 248731 209085 263877 209113
rect 263905 209085 263939 209113
rect 263967 209085 264001 209113
rect 264029 209085 264063 209113
rect 264091 209085 279237 209113
rect 279265 209085 279299 209113
rect 279327 209085 279361 209113
rect 279389 209085 279423 209113
rect 279451 209085 294597 209113
rect 294625 209085 294659 209113
rect 294687 209085 294721 209113
rect 294749 209085 294783 209113
rect 294811 209085 298248 209113
rect 298276 209085 298310 209113
rect 298338 209085 298372 209113
rect 298400 209085 298434 209113
rect 298462 209085 298990 209113
rect -958 209051 298990 209085
rect -958 209023 -430 209051
rect -402 209023 -368 209051
rect -340 209023 -306 209051
rect -278 209023 -244 209051
rect -216 209023 2757 209051
rect 2785 209023 2819 209051
rect 2847 209023 2881 209051
rect 2909 209023 2943 209051
rect 2971 209023 18117 209051
rect 18145 209023 18179 209051
rect 18207 209023 18241 209051
rect 18269 209023 18303 209051
rect 18331 209023 22259 209051
rect 22287 209023 22321 209051
rect 22349 209023 37619 209051
rect 37647 209023 37681 209051
rect 37709 209023 52979 209051
rect 53007 209023 53041 209051
rect 53069 209023 68339 209051
rect 68367 209023 68401 209051
rect 68429 209023 83699 209051
rect 83727 209023 83761 209051
rect 83789 209023 94917 209051
rect 94945 209023 94979 209051
rect 95007 209023 95041 209051
rect 95069 209023 95103 209051
rect 95131 209023 102259 209051
rect 102287 209023 102321 209051
rect 102349 209023 117619 209051
rect 117647 209023 117681 209051
rect 117709 209023 132979 209051
rect 133007 209023 133041 209051
rect 133069 209023 148339 209051
rect 148367 209023 148401 209051
rect 148429 209023 163699 209051
rect 163727 209023 163761 209051
rect 163789 209023 171717 209051
rect 171745 209023 171779 209051
rect 171807 209023 171841 209051
rect 171869 209023 171903 209051
rect 171931 209023 187077 209051
rect 187105 209023 187139 209051
rect 187167 209023 187201 209051
rect 187229 209023 187263 209051
rect 187291 209023 202437 209051
rect 202465 209023 202499 209051
rect 202527 209023 202561 209051
rect 202589 209023 202623 209051
rect 202651 209023 217797 209051
rect 217825 209023 217859 209051
rect 217887 209023 217921 209051
rect 217949 209023 217983 209051
rect 218011 209023 233157 209051
rect 233185 209023 233219 209051
rect 233247 209023 233281 209051
rect 233309 209023 233343 209051
rect 233371 209023 248517 209051
rect 248545 209023 248579 209051
rect 248607 209023 248641 209051
rect 248669 209023 248703 209051
rect 248731 209023 263877 209051
rect 263905 209023 263939 209051
rect 263967 209023 264001 209051
rect 264029 209023 264063 209051
rect 264091 209023 279237 209051
rect 279265 209023 279299 209051
rect 279327 209023 279361 209051
rect 279389 209023 279423 209051
rect 279451 209023 294597 209051
rect 294625 209023 294659 209051
rect 294687 209023 294721 209051
rect 294749 209023 294783 209051
rect 294811 209023 298248 209051
rect 298276 209023 298310 209051
rect 298338 209023 298372 209051
rect 298400 209023 298434 209051
rect 298462 209023 298990 209051
rect -958 208989 298990 209023
rect -958 208961 -430 208989
rect -402 208961 -368 208989
rect -340 208961 -306 208989
rect -278 208961 -244 208989
rect -216 208961 2757 208989
rect 2785 208961 2819 208989
rect 2847 208961 2881 208989
rect 2909 208961 2943 208989
rect 2971 208961 18117 208989
rect 18145 208961 18179 208989
rect 18207 208961 18241 208989
rect 18269 208961 18303 208989
rect 18331 208961 22259 208989
rect 22287 208961 22321 208989
rect 22349 208961 37619 208989
rect 37647 208961 37681 208989
rect 37709 208961 52979 208989
rect 53007 208961 53041 208989
rect 53069 208961 68339 208989
rect 68367 208961 68401 208989
rect 68429 208961 83699 208989
rect 83727 208961 83761 208989
rect 83789 208961 94917 208989
rect 94945 208961 94979 208989
rect 95007 208961 95041 208989
rect 95069 208961 95103 208989
rect 95131 208961 102259 208989
rect 102287 208961 102321 208989
rect 102349 208961 117619 208989
rect 117647 208961 117681 208989
rect 117709 208961 132979 208989
rect 133007 208961 133041 208989
rect 133069 208961 148339 208989
rect 148367 208961 148401 208989
rect 148429 208961 163699 208989
rect 163727 208961 163761 208989
rect 163789 208961 171717 208989
rect 171745 208961 171779 208989
rect 171807 208961 171841 208989
rect 171869 208961 171903 208989
rect 171931 208961 187077 208989
rect 187105 208961 187139 208989
rect 187167 208961 187201 208989
rect 187229 208961 187263 208989
rect 187291 208961 202437 208989
rect 202465 208961 202499 208989
rect 202527 208961 202561 208989
rect 202589 208961 202623 208989
rect 202651 208961 217797 208989
rect 217825 208961 217859 208989
rect 217887 208961 217921 208989
rect 217949 208961 217983 208989
rect 218011 208961 233157 208989
rect 233185 208961 233219 208989
rect 233247 208961 233281 208989
rect 233309 208961 233343 208989
rect 233371 208961 248517 208989
rect 248545 208961 248579 208989
rect 248607 208961 248641 208989
rect 248669 208961 248703 208989
rect 248731 208961 263877 208989
rect 263905 208961 263939 208989
rect 263967 208961 264001 208989
rect 264029 208961 264063 208989
rect 264091 208961 279237 208989
rect 279265 208961 279299 208989
rect 279327 208961 279361 208989
rect 279389 208961 279423 208989
rect 279451 208961 294597 208989
rect 294625 208961 294659 208989
rect 294687 208961 294721 208989
rect 294749 208961 294783 208989
rect 294811 208961 298248 208989
rect 298276 208961 298310 208989
rect 298338 208961 298372 208989
rect 298400 208961 298434 208989
rect 298462 208961 298990 208989
rect -958 208913 298990 208961
rect -958 203175 298990 203223
rect -958 203147 -910 203175
rect -882 203147 -848 203175
rect -820 203147 -786 203175
rect -758 203147 -724 203175
rect -696 203147 4617 203175
rect 4645 203147 4679 203175
rect 4707 203147 4741 203175
rect 4769 203147 4803 203175
rect 4831 203147 29939 203175
rect 29967 203147 30001 203175
rect 30029 203147 45299 203175
rect 45327 203147 45361 203175
rect 45389 203147 60659 203175
rect 60687 203147 60721 203175
rect 60749 203147 76019 203175
rect 76047 203147 76081 203175
rect 76109 203147 96777 203175
rect 96805 203147 96839 203175
rect 96867 203147 96901 203175
rect 96929 203147 96963 203175
rect 96991 203147 109939 203175
rect 109967 203147 110001 203175
rect 110029 203147 125299 203175
rect 125327 203147 125361 203175
rect 125389 203147 140659 203175
rect 140687 203147 140721 203175
rect 140749 203147 156019 203175
rect 156047 203147 156081 203175
rect 156109 203147 173577 203175
rect 173605 203147 173639 203175
rect 173667 203147 173701 203175
rect 173729 203147 173763 203175
rect 173791 203147 188937 203175
rect 188965 203147 188999 203175
rect 189027 203147 189061 203175
rect 189089 203147 189123 203175
rect 189151 203147 204297 203175
rect 204325 203147 204359 203175
rect 204387 203147 204421 203175
rect 204449 203147 204483 203175
rect 204511 203147 219657 203175
rect 219685 203147 219719 203175
rect 219747 203147 219781 203175
rect 219809 203147 219843 203175
rect 219871 203147 235017 203175
rect 235045 203147 235079 203175
rect 235107 203147 235141 203175
rect 235169 203147 235203 203175
rect 235231 203147 250377 203175
rect 250405 203147 250439 203175
rect 250467 203147 250501 203175
rect 250529 203147 250563 203175
rect 250591 203147 265737 203175
rect 265765 203147 265799 203175
rect 265827 203147 265861 203175
rect 265889 203147 265923 203175
rect 265951 203147 281097 203175
rect 281125 203147 281159 203175
rect 281187 203147 281221 203175
rect 281249 203147 281283 203175
rect 281311 203147 296457 203175
rect 296485 203147 296519 203175
rect 296547 203147 296581 203175
rect 296609 203147 296643 203175
rect 296671 203147 298728 203175
rect 298756 203147 298790 203175
rect 298818 203147 298852 203175
rect 298880 203147 298914 203175
rect 298942 203147 298990 203175
rect -958 203113 298990 203147
rect -958 203085 -910 203113
rect -882 203085 -848 203113
rect -820 203085 -786 203113
rect -758 203085 -724 203113
rect -696 203085 4617 203113
rect 4645 203085 4679 203113
rect 4707 203085 4741 203113
rect 4769 203085 4803 203113
rect 4831 203085 29939 203113
rect 29967 203085 30001 203113
rect 30029 203085 45299 203113
rect 45327 203085 45361 203113
rect 45389 203085 60659 203113
rect 60687 203085 60721 203113
rect 60749 203085 76019 203113
rect 76047 203085 76081 203113
rect 76109 203085 96777 203113
rect 96805 203085 96839 203113
rect 96867 203085 96901 203113
rect 96929 203085 96963 203113
rect 96991 203085 109939 203113
rect 109967 203085 110001 203113
rect 110029 203085 125299 203113
rect 125327 203085 125361 203113
rect 125389 203085 140659 203113
rect 140687 203085 140721 203113
rect 140749 203085 156019 203113
rect 156047 203085 156081 203113
rect 156109 203085 173577 203113
rect 173605 203085 173639 203113
rect 173667 203085 173701 203113
rect 173729 203085 173763 203113
rect 173791 203085 188937 203113
rect 188965 203085 188999 203113
rect 189027 203085 189061 203113
rect 189089 203085 189123 203113
rect 189151 203085 204297 203113
rect 204325 203085 204359 203113
rect 204387 203085 204421 203113
rect 204449 203085 204483 203113
rect 204511 203085 219657 203113
rect 219685 203085 219719 203113
rect 219747 203085 219781 203113
rect 219809 203085 219843 203113
rect 219871 203085 235017 203113
rect 235045 203085 235079 203113
rect 235107 203085 235141 203113
rect 235169 203085 235203 203113
rect 235231 203085 250377 203113
rect 250405 203085 250439 203113
rect 250467 203085 250501 203113
rect 250529 203085 250563 203113
rect 250591 203085 265737 203113
rect 265765 203085 265799 203113
rect 265827 203085 265861 203113
rect 265889 203085 265923 203113
rect 265951 203085 281097 203113
rect 281125 203085 281159 203113
rect 281187 203085 281221 203113
rect 281249 203085 281283 203113
rect 281311 203085 296457 203113
rect 296485 203085 296519 203113
rect 296547 203085 296581 203113
rect 296609 203085 296643 203113
rect 296671 203085 298728 203113
rect 298756 203085 298790 203113
rect 298818 203085 298852 203113
rect 298880 203085 298914 203113
rect 298942 203085 298990 203113
rect -958 203051 298990 203085
rect -958 203023 -910 203051
rect -882 203023 -848 203051
rect -820 203023 -786 203051
rect -758 203023 -724 203051
rect -696 203023 4617 203051
rect 4645 203023 4679 203051
rect 4707 203023 4741 203051
rect 4769 203023 4803 203051
rect 4831 203023 29939 203051
rect 29967 203023 30001 203051
rect 30029 203023 45299 203051
rect 45327 203023 45361 203051
rect 45389 203023 60659 203051
rect 60687 203023 60721 203051
rect 60749 203023 76019 203051
rect 76047 203023 76081 203051
rect 76109 203023 96777 203051
rect 96805 203023 96839 203051
rect 96867 203023 96901 203051
rect 96929 203023 96963 203051
rect 96991 203023 109939 203051
rect 109967 203023 110001 203051
rect 110029 203023 125299 203051
rect 125327 203023 125361 203051
rect 125389 203023 140659 203051
rect 140687 203023 140721 203051
rect 140749 203023 156019 203051
rect 156047 203023 156081 203051
rect 156109 203023 173577 203051
rect 173605 203023 173639 203051
rect 173667 203023 173701 203051
rect 173729 203023 173763 203051
rect 173791 203023 188937 203051
rect 188965 203023 188999 203051
rect 189027 203023 189061 203051
rect 189089 203023 189123 203051
rect 189151 203023 204297 203051
rect 204325 203023 204359 203051
rect 204387 203023 204421 203051
rect 204449 203023 204483 203051
rect 204511 203023 219657 203051
rect 219685 203023 219719 203051
rect 219747 203023 219781 203051
rect 219809 203023 219843 203051
rect 219871 203023 235017 203051
rect 235045 203023 235079 203051
rect 235107 203023 235141 203051
rect 235169 203023 235203 203051
rect 235231 203023 250377 203051
rect 250405 203023 250439 203051
rect 250467 203023 250501 203051
rect 250529 203023 250563 203051
rect 250591 203023 265737 203051
rect 265765 203023 265799 203051
rect 265827 203023 265861 203051
rect 265889 203023 265923 203051
rect 265951 203023 281097 203051
rect 281125 203023 281159 203051
rect 281187 203023 281221 203051
rect 281249 203023 281283 203051
rect 281311 203023 296457 203051
rect 296485 203023 296519 203051
rect 296547 203023 296581 203051
rect 296609 203023 296643 203051
rect 296671 203023 298728 203051
rect 298756 203023 298790 203051
rect 298818 203023 298852 203051
rect 298880 203023 298914 203051
rect 298942 203023 298990 203051
rect -958 202989 298990 203023
rect -958 202961 -910 202989
rect -882 202961 -848 202989
rect -820 202961 -786 202989
rect -758 202961 -724 202989
rect -696 202961 4617 202989
rect 4645 202961 4679 202989
rect 4707 202961 4741 202989
rect 4769 202961 4803 202989
rect 4831 202961 29939 202989
rect 29967 202961 30001 202989
rect 30029 202961 45299 202989
rect 45327 202961 45361 202989
rect 45389 202961 60659 202989
rect 60687 202961 60721 202989
rect 60749 202961 76019 202989
rect 76047 202961 76081 202989
rect 76109 202961 96777 202989
rect 96805 202961 96839 202989
rect 96867 202961 96901 202989
rect 96929 202961 96963 202989
rect 96991 202961 109939 202989
rect 109967 202961 110001 202989
rect 110029 202961 125299 202989
rect 125327 202961 125361 202989
rect 125389 202961 140659 202989
rect 140687 202961 140721 202989
rect 140749 202961 156019 202989
rect 156047 202961 156081 202989
rect 156109 202961 173577 202989
rect 173605 202961 173639 202989
rect 173667 202961 173701 202989
rect 173729 202961 173763 202989
rect 173791 202961 188937 202989
rect 188965 202961 188999 202989
rect 189027 202961 189061 202989
rect 189089 202961 189123 202989
rect 189151 202961 204297 202989
rect 204325 202961 204359 202989
rect 204387 202961 204421 202989
rect 204449 202961 204483 202989
rect 204511 202961 219657 202989
rect 219685 202961 219719 202989
rect 219747 202961 219781 202989
rect 219809 202961 219843 202989
rect 219871 202961 235017 202989
rect 235045 202961 235079 202989
rect 235107 202961 235141 202989
rect 235169 202961 235203 202989
rect 235231 202961 250377 202989
rect 250405 202961 250439 202989
rect 250467 202961 250501 202989
rect 250529 202961 250563 202989
rect 250591 202961 265737 202989
rect 265765 202961 265799 202989
rect 265827 202961 265861 202989
rect 265889 202961 265923 202989
rect 265951 202961 281097 202989
rect 281125 202961 281159 202989
rect 281187 202961 281221 202989
rect 281249 202961 281283 202989
rect 281311 202961 296457 202989
rect 296485 202961 296519 202989
rect 296547 202961 296581 202989
rect 296609 202961 296643 202989
rect 296671 202961 298728 202989
rect 298756 202961 298790 202989
rect 298818 202961 298852 202989
rect 298880 202961 298914 202989
rect 298942 202961 298990 202989
rect -958 202913 298990 202961
rect -958 200175 298990 200223
rect -958 200147 -430 200175
rect -402 200147 -368 200175
rect -340 200147 -306 200175
rect -278 200147 -244 200175
rect -216 200147 2757 200175
rect 2785 200147 2819 200175
rect 2847 200147 2881 200175
rect 2909 200147 2943 200175
rect 2971 200147 18117 200175
rect 18145 200147 18179 200175
rect 18207 200147 18241 200175
rect 18269 200147 18303 200175
rect 18331 200147 22259 200175
rect 22287 200147 22321 200175
rect 22349 200147 37619 200175
rect 37647 200147 37681 200175
rect 37709 200147 52979 200175
rect 53007 200147 53041 200175
rect 53069 200147 68339 200175
rect 68367 200147 68401 200175
rect 68429 200147 83699 200175
rect 83727 200147 83761 200175
rect 83789 200147 94917 200175
rect 94945 200147 94979 200175
rect 95007 200147 95041 200175
rect 95069 200147 95103 200175
rect 95131 200147 102259 200175
rect 102287 200147 102321 200175
rect 102349 200147 117619 200175
rect 117647 200147 117681 200175
rect 117709 200147 132979 200175
rect 133007 200147 133041 200175
rect 133069 200147 148339 200175
rect 148367 200147 148401 200175
rect 148429 200147 163699 200175
rect 163727 200147 163761 200175
rect 163789 200147 171717 200175
rect 171745 200147 171779 200175
rect 171807 200147 171841 200175
rect 171869 200147 171903 200175
rect 171931 200147 187077 200175
rect 187105 200147 187139 200175
rect 187167 200147 187201 200175
rect 187229 200147 187263 200175
rect 187291 200147 202437 200175
rect 202465 200147 202499 200175
rect 202527 200147 202561 200175
rect 202589 200147 202623 200175
rect 202651 200147 217797 200175
rect 217825 200147 217859 200175
rect 217887 200147 217921 200175
rect 217949 200147 217983 200175
rect 218011 200147 233157 200175
rect 233185 200147 233219 200175
rect 233247 200147 233281 200175
rect 233309 200147 233343 200175
rect 233371 200147 248517 200175
rect 248545 200147 248579 200175
rect 248607 200147 248641 200175
rect 248669 200147 248703 200175
rect 248731 200147 263877 200175
rect 263905 200147 263939 200175
rect 263967 200147 264001 200175
rect 264029 200147 264063 200175
rect 264091 200147 279237 200175
rect 279265 200147 279299 200175
rect 279327 200147 279361 200175
rect 279389 200147 279423 200175
rect 279451 200147 294597 200175
rect 294625 200147 294659 200175
rect 294687 200147 294721 200175
rect 294749 200147 294783 200175
rect 294811 200147 298248 200175
rect 298276 200147 298310 200175
rect 298338 200147 298372 200175
rect 298400 200147 298434 200175
rect 298462 200147 298990 200175
rect -958 200113 298990 200147
rect -958 200085 -430 200113
rect -402 200085 -368 200113
rect -340 200085 -306 200113
rect -278 200085 -244 200113
rect -216 200085 2757 200113
rect 2785 200085 2819 200113
rect 2847 200085 2881 200113
rect 2909 200085 2943 200113
rect 2971 200085 18117 200113
rect 18145 200085 18179 200113
rect 18207 200085 18241 200113
rect 18269 200085 18303 200113
rect 18331 200085 22259 200113
rect 22287 200085 22321 200113
rect 22349 200085 37619 200113
rect 37647 200085 37681 200113
rect 37709 200085 52979 200113
rect 53007 200085 53041 200113
rect 53069 200085 68339 200113
rect 68367 200085 68401 200113
rect 68429 200085 83699 200113
rect 83727 200085 83761 200113
rect 83789 200085 94917 200113
rect 94945 200085 94979 200113
rect 95007 200085 95041 200113
rect 95069 200085 95103 200113
rect 95131 200085 102259 200113
rect 102287 200085 102321 200113
rect 102349 200085 117619 200113
rect 117647 200085 117681 200113
rect 117709 200085 132979 200113
rect 133007 200085 133041 200113
rect 133069 200085 148339 200113
rect 148367 200085 148401 200113
rect 148429 200085 163699 200113
rect 163727 200085 163761 200113
rect 163789 200085 171717 200113
rect 171745 200085 171779 200113
rect 171807 200085 171841 200113
rect 171869 200085 171903 200113
rect 171931 200085 187077 200113
rect 187105 200085 187139 200113
rect 187167 200085 187201 200113
rect 187229 200085 187263 200113
rect 187291 200085 202437 200113
rect 202465 200085 202499 200113
rect 202527 200085 202561 200113
rect 202589 200085 202623 200113
rect 202651 200085 217797 200113
rect 217825 200085 217859 200113
rect 217887 200085 217921 200113
rect 217949 200085 217983 200113
rect 218011 200085 233157 200113
rect 233185 200085 233219 200113
rect 233247 200085 233281 200113
rect 233309 200085 233343 200113
rect 233371 200085 248517 200113
rect 248545 200085 248579 200113
rect 248607 200085 248641 200113
rect 248669 200085 248703 200113
rect 248731 200085 263877 200113
rect 263905 200085 263939 200113
rect 263967 200085 264001 200113
rect 264029 200085 264063 200113
rect 264091 200085 279237 200113
rect 279265 200085 279299 200113
rect 279327 200085 279361 200113
rect 279389 200085 279423 200113
rect 279451 200085 294597 200113
rect 294625 200085 294659 200113
rect 294687 200085 294721 200113
rect 294749 200085 294783 200113
rect 294811 200085 298248 200113
rect 298276 200085 298310 200113
rect 298338 200085 298372 200113
rect 298400 200085 298434 200113
rect 298462 200085 298990 200113
rect -958 200051 298990 200085
rect -958 200023 -430 200051
rect -402 200023 -368 200051
rect -340 200023 -306 200051
rect -278 200023 -244 200051
rect -216 200023 2757 200051
rect 2785 200023 2819 200051
rect 2847 200023 2881 200051
rect 2909 200023 2943 200051
rect 2971 200023 18117 200051
rect 18145 200023 18179 200051
rect 18207 200023 18241 200051
rect 18269 200023 18303 200051
rect 18331 200023 22259 200051
rect 22287 200023 22321 200051
rect 22349 200023 37619 200051
rect 37647 200023 37681 200051
rect 37709 200023 52979 200051
rect 53007 200023 53041 200051
rect 53069 200023 68339 200051
rect 68367 200023 68401 200051
rect 68429 200023 83699 200051
rect 83727 200023 83761 200051
rect 83789 200023 94917 200051
rect 94945 200023 94979 200051
rect 95007 200023 95041 200051
rect 95069 200023 95103 200051
rect 95131 200023 102259 200051
rect 102287 200023 102321 200051
rect 102349 200023 117619 200051
rect 117647 200023 117681 200051
rect 117709 200023 132979 200051
rect 133007 200023 133041 200051
rect 133069 200023 148339 200051
rect 148367 200023 148401 200051
rect 148429 200023 163699 200051
rect 163727 200023 163761 200051
rect 163789 200023 171717 200051
rect 171745 200023 171779 200051
rect 171807 200023 171841 200051
rect 171869 200023 171903 200051
rect 171931 200023 187077 200051
rect 187105 200023 187139 200051
rect 187167 200023 187201 200051
rect 187229 200023 187263 200051
rect 187291 200023 202437 200051
rect 202465 200023 202499 200051
rect 202527 200023 202561 200051
rect 202589 200023 202623 200051
rect 202651 200023 217797 200051
rect 217825 200023 217859 200051
rect 217887 200023 217921 200051
rect 217949 200023 217983 200051
rect 218011 200023 233157 200051
rect 233185 200023 233219 200051
rect 233247 200023 233281 200051
rect 233309 200023 233343 200051
rect 233371 200023 248517 200051
rect 248545 200023 248579 200051
rect 248607 200023 248641 200051
rect 248669 200023 248703 200051
rect 248731 200023 263877 200051
rect 263905 200023 263939 200051
rect 263967 200023 264001 200051
rect 264029 200023 264063 200051
rect 264091 200023 279237 200051
rect 279265 200023 279299 200051
rect 279327 200023 279361 200051
rect 279389 200023 279423 200051
rect 279451 200023 294597 200051
rect 294625 200023 294659 200051
rect 294687 200023 294721 200051
rect 294749 200023 294783 200051
rect 294811 200023 298248 200051
rect 298276 200023 298310 200051
rect 298338 200023 298372 200051
rect 298400 200023 298434 200051
rect 298462 200023 298990 200051
rect -958 199989 298990 200023
rect -958 199961 -430 199989
rect -402 199961 -368 199989
rect -340 199961 -306 199989
rect -278 199961 -244 199989
rect -216 199961 2757 199989
rect 2785 199961 2819 199989
rect 2847 199961 2881 199989
rect 2909 199961 2943 199989
rect 2971 199961 18117 199989
rect 18145 199961 18179 199989
rect 18207 199961 18241 199989
rect 18269 199961 18303 199989
rect 18331 199961 22259 199989
rect 22287 199961 22321 199989
rect 22349 199961 37619 199989
rect 37647 199961 37681 199989
rect 37709 199961 52979 199989
rect 53007 199961 53041 199989
rect 53069 199961 68339 199989
rect 68367 199961 68401 199989
rect 68429 199961 83699 199989
rect 83727 199961 83761 199989
rect 83789 199961 94917 199989
rect 94945 199961 94979 199989
rect 95007 199961 95041 199989
rect 95069 199961 95103 199989
rect 95131 199961 102259 199989
rect 102287 199961 102321 199989
rect 102349 199961 117619 199989
rect 117647 199961 117681 199989
rect 117709 199961 132979 199989
rect 133007 199961 133041 199989
rect 133069 199961 148339 199989
rect 148367 199961 148401 199989
rect 148429 199961 163699 199989
rect 163727 199961 163761 199989
rect 163789 199961 171717 199989
rect 171745 199961 171779 199989
rect 171807 199961 171841 199989
rect 171869 199961 171903 199989
rect 171931 199961 187077 199989
rect 187105 199961 187139 199989
rect 187167 199961 187201 199989
rect 187229 199961 187263 199989
rect 187291 199961 202437 199989
rect 202465 199961 202499 199989
rect 202527 199961 202561 199989
rect 202589 199961 202623 199989
rect 202651 199961 217797 199989
rect 217825 199961 217859 199989
rect 217887 199961 217921 199989
rect 217949 199961 217983 199989
rect 218011 199961 233157 199989
rect 233185 199961 233219 199989
rect 233247 199961 233281 199989
rect 233309 199961 233343 199989
rect 233371 199961 248517 199989
rect 248545 199961 248579 199989
rect 248607 199961 248641 199989
rect 248669 199961 248703 199989
rect 248731 199961 263877 199989
rect 263905 199961 263939 199989
rect 263967 199961 264001 199989
rect 264029 199961 264063 199989
rect 264091 199961 279237 199989
rect 279265 199961 279299 199989
rect 279327 199961 279361 199989
rect 279389 199961 279423 199989
rect 279451 199961 294597 199989
rect 294625 199961 294659 199989
rect 294687 199961 294721 199989
rect 294749 199961 294783 199989
rect 294811 199961 298248 199989
rect 298276 199961 298310 199989
rect 298338 199961 298372 199989
rect 298400 199961 298434 199989
rect 298462 199961 298990 199989
rect -958 199913 298990 199961
rect -958 194175 298990 194223
rect -958 194147 -910 194175
rect -882 194147 -848 194175
rect -820 194147 -786 194175
rect -758 194147 -724 194175
rect -696 194147 4617 194175
rect 4645 194147 4679 194175
rect 4707 194147 4741 194175
rect 4769 194147 4803 194175
rect 4831 194147 29939 194175
rect 29967 194147 30001 194175
rect 30029 194147 45299 194175
rect 45327 194147 45361 194175
rect 45389 194147 60659 194175
rect 60687 194147 60721 194175
rect 60749 194147 76019 194175
rect 76047 194147 76081 194175
rect 76109 194147 96777 194175
rect 96805 194147 96839 194175
rect 96867 194147 96901 194175
rect 96929 194147 96963 194175
rect 96991 194147 109939 194175
rect 109967 194147 110001 194175
rect 110029 194147 125299 194175
rect 125327 194147 125361 194175
rect 125389 194147 140659 194175
rect 140687 194147 140721 194175
rect 140749 194147 156019 194175
rect 156047 194147 156081 194175
rect 156109 194147 173577 194175
rect 173605 194147 173639 194175
rect 173667 194147 173701 194175
rect 173729 194147 173763 194175
rect 173791 194147 188937 194175
rect 188965 194147 188999 194175
rect 189027 194147 189061 194175
rect 189089 194147 189123 194175
rect 189151 194147 189939 194175
rect 189967 194147 190001 194175
rect 190029 194147 204297 194175
rect 204325 194147 204359 194175
rect 204387 194147 204421 194175
rect 204449 194147 204483 194175
rect 204511 194147 219657 194175
rect 219685 194147 219719 194175
rect 219747 194147 219781 194175
rect 219809 194147 219843 194175
rect 219871 194147 235017 194175
rect 235045 194147 235079 194175
rect 235107 194147 235141 194175
rect 235169 194147 235203 194175
rect 235231 194147 250377 194175
rect 250405 194147 250439 194175
rect 250467 194147 250501 194175
rect 250529 194147 250563 194175
rect 250591 194147 265737 194175
rect 265765 194147 265799 194175
rect 265827 194147 265861 194175
rect 265889 194147 265923 194175
rect 265951 194147 281097 194175
rect 281125 194147 281159 194175
rect 281187 194147 281221 194175
rect 281249 194147 281283 194175
rect 281311 194147 296457 194175
rect 296485 194147 296519 194175
rect 296547 194147 296581 194175
rect 296609 194147 296643 194175
rect 296671 194147 298728 194175
rect 298756 194147 298790 194175
rect 298818 194147 298852 194175
rect 298880 194147 298914 194175
rect 298942 194147 298990 194175
rect -958 194113 298990 194147
rect -958 194085 -910 194113
rect -882 194085 -848 194113
rect -820 194085 -786 194113
rect -758 194085 -724 194113
rect -696 194085 4617 194113
rect 4645 194085 4679 194113
rect 4707 194085 4741 194113
rect 4769 194085 4803 194113
rect 4831 194085 29939 194113
rect 29967 194085 30001 194113
rect 30029 194085 45299 194113
rect 45327 194085 45361 194113
rect 45389 194085 60659 194113
rect 60687 194085 60721 194113
rect 60749 194085 76019 194113
rect 76047 194085 76081 194113
rect 76109 194085 96777 194113
rect 96805 194085 96839 194113
rect 96867 194085 96901 194113
rect 96929 194085 96963 194113
rect 96991 194085 109939 194113
rect 109967 194085 110001 194113
rect 110029 194085 125299 194113
rect 125327 194085 125361 194113
rect 125389 194085 140659 194113
rect 140687 194085 140721 194113
rect 140749 194085 156019 194113
rect 156047 194085 156081 194113
rect 156109 194085 173577 194113
rect 173605 194085 173639 194113
rect 173667 194085 173701 194113
rect 173729 194085 173763 194113
rect 173791 194085 188937 194113
rect 188965 194085 188999 194113
rect 189027 194085 189061 194113
rect 189089 194085 189123 194113
rect 189151 194085 189939 194113
rect 189967 194085 190001 194113
rect 190029 194085 204297 194113
rect 204325 194085 204359 194113
rect 204387 194085 204421 194113
rect 204449 194085 204483 194113
rect 204511 194085 219657 194113
rect 219685 194085 219719 194113
rect 219747 194085 219781 194113
rect 219809 194085 219843 194113
rect 219871 194085 235017 194113
rect 235045 194085 235079 194113
rect 235107 194085 235141 194113
rect 235169 194085 235203 194113
rect 235231 194085 250377 194113
rect 250405 194085 250439 194113
rect 250467 194085 250501 194113
rect 250529 194085 250563 194113
rect 250591 194085 265737 194113
rect 265765 194085 265799 194113
rect 265827 194085 265861 194113
rect 265889 194085 265923 194113
rect 265951 194085 281097 194113
rect 281125 194085 281159 194113
rect 281187 194085 281221 194113
rect 281249 194085 281283 194113
rect 281311 194085 296457 194113
rect 296485 194085 296519 194113
rect 296547 194085 296581 194113
rect 296609 194085 296643 194113
rect 296671 194085 298728 194113
rect 298756 194085 298790 194113
rect 298818 194085 298852 194113
rect 298880 194085 298914 194113
rect 298942 194085 298990 194113
rect -958 194051 298990 194085
rect -958 194023 -910 194051
rect -882 194023 -848 194051
rect -820 194023 -786 194051
rect -758 194023 -724 194051
rect -696 194023 4617 194051
rect 4645 194023 4679 194051
rect 4707 194023 4741 194051
rect 4769 194023 4803 194051
rect 4831 194023 29939 194051
rect 29967 194023 30001 194051
rect 30029 194023 45299 194051
rect 45327 194023 45361 194051
rect 45389 194023 60659 194051
rect 60687 194023 60721 194051
rect 60749 194023 76019 194051
rect 76047 194023 76081 194051
rect 76109 194023 96777 194051
rect 96805 194023 96839 194051
rect 96867 194023 96901 194051
rect 96929 194023 96963 194051
rect 96991 194023 109939 194051
rect 109967 194023 110001 194051
rect 110029 194023 125299 194051
rect 125327 194023 125361 194051
rect 125389 194023 140659 194051
rect 140687 194023 140721 194051
rect 140749 194023 156019 194051
rect 156047 194023 156081 194051
rect 156109 194023 173577 194051
rect 173605 194023 173639 194051
rect 173667 194023 173701 194051
rect 173729 194023 173763 194051
rect 173791 194023 188937 194051
rect 188965 194023 188999 194051
rect 189027 194023 189061 194051
rect 189089 194023 189123 194051
rect 189151 194023 189939 194051
rect 189967 194023 190001 194051
rect 190029 194023 204297 194051
rect 204325 194023 204359 194051
rect 204387 194023 204421 194051
rect 204449 194023 204483 194051
rect 204511 194023 219657 194051
rect 219685 194023 219719 194051
rect 219747 194023 219781 194051
rect 219809 194023 219843 194051
rect 219871 194023 235017 194051
rect 235045 194023 235079 194051
rect 235107 194023 235141 194051
rect 235169 194023 235203 194051
rect 235231 194023 250377 194051
rect 250405 194023 250439 194051
rect 250467 194023 250501 194051
rect 250529 194023 250563 194051
rect 250591 194023 265737 194051
rect 265765 194023 265799 194051
rect 265827 194023 265861 194051
rect 265889 194023 265923 194051
rect 265951 194023 281097 194051
rect 281125 194023 281159 194051
rect 281187 194023 281221 194051
rect 281249 194023 281283 194051
rect 281311 194023 296457 194051
rect 296485 194023 296519 194051
rect 296547 194023 296581 194051
rect 296609 194023 296643 194051
rect 296671 194023 298728 194051
rect 298756 194023 298790 194051
rect 298818 194023 298852 194051
rect 298880 194023 298914 194051
rect 298942 194023 298990 194051
rect -958 193989 298990 194023
rect -958 193961 -910 193989
rect -882 193961 -848 193989
rect -820 193961 -786 193989
rect -758 193961 -724 193989
rect -696 193961 4617 193989
rect 4645 193961 4679 193989
rect 4707 193961 4741 193989
rect 4769 193961 4803 193989
rect 4831 193961 29939 193989
rect 29967 193961 30001 193989
rect 30029 193961 45299 193989
rect 45327 193961 45361 193989
rect 45389 193961 60659 193989
rect 60687 193961 60721 193989
rect 60749 193961 76019 193989
rect 76047 193961 76081 193989
rect 76109 193961 96777 193989
rect 96805 193961 96839 193989
rect 96867 193961 96901 193989
rect 96929 193961 96963 193989
rect 96991 193961 109939 193989
rect 109967 193961 110001 193989
rect 110029 193961 125299 193989
rect 125327 193961 125361 193989
rect 125389 193961 140659 193989
rect 140687 193961 140721 193989
rect 140749 193961 156019 193989
rect 156047 193961 156081 193989
rect 156109 193961 173577 193989
rect 173605 193961 173639 193989
rect 173667 193961 173701 193989
rect 173729 193961 173763 193989
rect 173791 193961 188937 193989
rect 188965 193961 188999 193989
rect 189027 193961 189061 193989
rect 189089 193961 189123 193989
rect 189151 193961 189939 193989
rect 189967 193961 190001 193989
rect 190029 193961 204297 193989
rect 204325 193961 204359 193989
rect 204387 193961 204421 193989
rect 204449 193961 204483 193989
rect 204511 193961 219657 193989
rect 219685 193961 219719 193989
rect 219747 193961 219781 193989
rect 219809 193961 219843 193989
rect 219871 193961 235017 193989
rect 235045 193961 235079 193989
rect 235107 193961 235141 193989
rect 235169 193961 235203 193989
rect 235231 193961 250377 193989
rect 250405 193961 250439 193989
rect 250467 193961 250501 193989
rect 250529 193961 250563 193989
rect 250591 193961 265737 193989
rect 265765 193961 265799 193989
rect 265827 193961 265861 193989
rect 265889 193961 265923 193989
rect 265951 193961 281097 193989
rect 281125 193961 281159 193989
rect 281187 193961 281221 193989
rect 281249 193961 281283 193989
rect 281311 193961 296457 193989
rect 296485 193961 296519 193989
rect 296547 193961 296581 193989
rect 296609 193961 296643 193989
rect 296671 193961 298728 193989
rect 298756 193961 298790 193989
rect 298818 193961 298852 193989
rect 298880 193961 298914 193989
rect 298942 193961 298990 193989
rect -958 193913 298990 193961
rect -958 191175 298990 191223
rect -958 191147 -430 191175
rect -402 191147 -368 191175
rect -340 191147 -306 191175
rect -278 191147 -244 191175
rect -216 191147 2757 191175
rect 2785 191147 2819 191175
rect 2847 191147 2881 191175
rect 2909 191147 2943 191175
rect 2971 191147 18117 191175
rect 18145 191147 18179 191175
rect 18207 191147 18241 191175
rect 18269 191147 18303 191175
rect 18331 191147 22259 191175
rect 22287 191147 22321 191175
rect 22349 191147 37619 191175
rect 37647 191147 37681 191175
rect 37709 191147 52979 191175
rect 53007 191147 53041 191175
rect 53069 191147 68339 191175
rect 68367 191147 68401 191175
rect 68429 191147 83699 191175
rect 83727 191147 83761 191175
rect 83789 191147 94917 191175
rect 94945 191147 94979 191175
rect 95007 191147 95041 191175
rect 95069 191147 95103 191175
rect 95131 191147 102259 191175
rect 102287 191147 102321 191175
rect 102349 191147 117619 191175
rect 117647 191147 117681 191175
rect 117709 191147 132979 191175
rect 133007 191147 133041 191175
rect 133069 191147 148339 191175
rect 148367 191147 148401 191175
rect 148429 191147 163699 191175
rect 163727 191147 163761 191175
rect 163789 191147 171717 191175
rect 171745 191147 171779 191175
rect 171807 191147 171841 191175
rect 171869 191147 171903 191175
rect 171931 191147 182259 191175
rect 182287 191147 182321 191175
rect 182349 191147 197619 191175
rect 197647 191147 197681 191175
rect 197709 191147 202437 191175
rect 202465 191147 202499 191175
rect 202527 191147 202561 191175
rect 202589 191147 202623 191175
rect 202651 191147 217797 191175
rect 217825 191147 217859 191175
rect 217887 191147 217921 191175
rect 217949 191147 217983 191175
rect 218011 191147 233157 191175
rect 233185 191147 233219 191175
rect 233247 191147 233281 191175
rect 233309 191147 233343 191175
rect 233371 191147 248517 191175
rect 248545 191147 248579 191175
rect 248607 191147 248641 191175
rect 248669 191147 248703 191175
rect 248731 191147 263877 191175
rect 263905 191147 263939 191175
rect 263967 191147 264001 191175
rect 264029 191147 264063 191175
rect 264091 191147 279237 191175
rect 279265 191147 279299 191175
rect 279327 191147 279361 191175
rect 279389 191147 279423 191175
rect 279451 191147 294597 191175
rect 294625 191147 294659 191175
rect 294687 191147 294721 191175
rect 294749 191147 294783 191175
rect 294811 191147 298248 191175
rect 298276 191147 298310 191175
rect 298338 191147 298372 191175
rect 298400 191147 298434 191175
rect 298462 191147 298990 191175
rect -958 191113 298990 191147
rect -958 191085 -430 191113
rect -402 191085 -368 191113
rect -340 191085 -306 191113
rect -278 191085 -244 191113
rect -216 191085 2757 191113
rect 2785 191085 2819 191113
rect 2847 191085 2881 191113
rect 2909 191085 2943 191113
rect 2971 191085 18117 191113
rect 18145 191085 18179 191113
rect 18207 191085 18241 191113
rect 18269 191085 18303 191113
rect 18331 191085 22259 191113
rect 22287 191085 22321 191113
rect 22349 191085 37619 191113
rect 37647 191085 37681 191113
rect 37709 191085 52979 191113
rect 53007 191085 53041 191113
rect 53069 191085 68339 191113
rect 68367 191085 68401 191113
rect 68429 191085 83699 191113
rect 83727 191085 83761 191113
rect 83789 191085 94917 191113
rect 94945 191085 94979 191113
rect 95007 191085 95041 191113
rect 95069 191085 95103 191113
rect 95131 191085 102259 191113
rect 102287 191085 102321 191113
rect 102349 191085 117619 191113
rect 117647 191085 117681 191113
rect 117709 191085 132979 191113
rect 133007 191085 133041 191113
rect 133069 191085 148339 191113
rect 148367 191085 148401 191113
rect 148429 191085 163699 191113
rect 163727 191085 163761 191113
rect 163789 191085 171717 191113
rect 171745 191085 171779 191113
rect 171807 191085 171841 191113
rect 171869 191085 171903 191113
rect 171931 191085 182259 191113
rect 182287 191085 182321 191113
rect 182349 191085 197619 191113
rect 197647 191085 197681 191113
rect 197709 191085 202437 191113
rect 202465 191085 202499 191113
rect 202527 191085 202561 191113
rect 202589 191085 202623 191113
rect 202651 191085 217797 191113
rect 217825 191085 217859 191113
rect 217887 191085 217921 191113
rect 217949 191085 217983 191113
rect 218011 191085 233157 191113
rect 233185 191085 233219 191113
rect 233247 191085 233281 191113
rect 233309 191085 233343 191113
rect 233371 191085 248517 191113
rect 248545 191085 248579 191113
rect 248607 191085 248641 191113
rect 248669 191085 248703 191113
rect 248731 191085 263877 191113
rect 263905 191085 263939 191113
rect 263967 191085 264001 191113
rect 264029 191085 264063 191113
rect 264091 191085 279237 191113
rect 279265 191085 279299 191113
rect 279327 191085 279361 191113
rect 279389 191085 279423 191113
rect 279451 191085 294597 191113
rect 294625 191085 294659 191113
rect 294687 191085 294721 191113
rect 294749 191085 294783 191113
rect 294811 191085 298248 191113
rect 298276 191085 298310 191113
rect 298338 191085 298372 191113
rect 298400 191085 298434 191113
rect 298462 191085 298990 191113
rect -958 191051 298990 191085
rect -958 191023 -430 191051
rect -402 191023 -368 191051
rect -340 191023 -306 191051
rect -278 191023 -244 191051
rect -216 191023 2757 191051
rect 2785 191023 2819 191051
rect 2847 191023 2881 191051
rect 2909 191023 2943 191051
rect 2971 191023 18117 191051
rect 18145 191023 18179 191051
rect 18207 191023 18241 191051
rect 18269 191023 18303 191051
rect 18331 191023 22259 191051
rect 22287 191023 22321 191051
rect 22349 191023 37619 191051
rect 37647 191023 37681 191051
rect 37709 191023 52979 191051
rect 53007 191023 53041 191051
rect 53069 191023 68339 191051
rect 68367 191023 68401 191051
rect 68429 191023 83699 191051
rect 83727 191023 83761 191051
rect 83789 191023 94917 191051
rect 94945 191023 94979 191051
rect 95007 191023 95041 191051
rect 95069 191023 95103 191051
rect 95131 191023 102259 191051
rect 102287 191023 102321 191051
rect 102349 191023 117619 191051
rect 117647 191023 117681 191051
rect 117709 191023 132979 191051
rect 133007 191023 133041 191051
rect 133069 191023 148339 191051
rect 148367 191023 148401 191051
rect 148429 191023 163699 191051
rect 163727 191023 163761 191051
rect 163789 191023 171717 191051
rect 171745 191023 171779 191051
rect 171807 191023 171841 191051
rect 171869 191023 171903 191051
rect 171931 191023 182259 191051
rect 182287 191023 182321 191051
rect 182349 191023 197619 191051
rect 197647 191023 197681 191051
rect 197709 191023 202437 191051
rect 202465 191023 202499 191051
rect 202527 191023 202561 191051
rect 202589 191023 202623 191051
rect 202651 191023 217797 191051
rect 217825 191023 217859 191051
rect 217887 191023 217921 191051
rect 217949 191023 217983 191051
rect 218011 191023 233157 191051
rect 233185 191023 233219 191051
rect 233247 191023 233281 191051
rect 233309 191023 233343 191051
rect 233371 191023 248517 191051
rect 248545 191023 248579 191051
rect 248607 191023 248641 191051
rect 248669 191023 248703 191051
rect 248731 191023 263877 191051
rect 263905 191023 263939 191051
rect 263967 191023 264001 191051
rect 264029 191023 264063 191051
rect 264091 191023 279237 191051
rect 279265 191023 279299 191051
rect 279327 191023 279361 191051
rect 279389 191023 279423 191051
rect 279451 191023 294597 191051
rect 294625 191023 294659 191051
rect 294687 191023 294721 191051
rect 294749 191023 294783 191051
rect 294811 191023 298248 191051
rect 298276 191023 298310 191051
rect 298338 191023 298372 191051
rect 298400 191023 298434 191051
rect 298462 191023 298990 191051
rect -958 190989 298990 191023
rect -958 190961 -430 190989
rect -402 190961 -368 190989
rect -340 190961 -306 190989
rect -278 190961 -244 190989
rect -216 190961 2757 190989
rect 2785 190961 2819 190989
rect 2847 190961 2881 190989
rect 2909 190961 2943 190989
rect 2971 190961 18117 190989
rect 18145 190961 18179 190989
rect 18207 190961 18241 190989
rect 18269 190961 18303 190989
rect 18331 190961 22259 190989
rect 22287 190961 22321 190989
rect 22349 190961 37619 190989
rect 37647 190961 37681 190989
rect 37709 190961 52979 190989
rect 53007 190961 53041 190989
rect 53069 190961 68339 190989
rect 68367 190961 68401 190989
rect 68429 190961 83699 190989
rect 83727 190961 83761 190989
rect 83789 190961 94917 190989
rect 94945 190961 94979 190989
rect 95007 190961 95041 190989
rect 95069 190961 95103 190989
rect 95131 190961 102259 190989
rect 102287 190961 102321 190989
rect 102349 190961 117619 190989
rect 117647 190961 117681 190989
rect 117709 190961 132979 190989
rect 133007 190961 133041 190989
rect 133069 190961 148339 190989
rect 148367 190961 148401 190989
rect 148429 190961 163699 190989
rect 163727 190961 163761 190989
rect 163789 190961 171717 190989
rect 171745 190961 171779 190989
rect 171807 190961 171841 190989
rect 171869 190961 171903 190989
rect 171931 190961 182259 190989
rect 182287 190961 182321 190989
rect 182349 190961 197619 190989
rect 197647 190961 197681 190989
rect 197709 190961 202437 190989
rect 202465 190961 202499 190989
rect 202527 190961 202561 190989
rect 202589 190961 202623 190989
rect 202651 190961 217797 190989
rect 217825 190961 217859 190989
rect 217887 190961 217921 190989
rect 217949 190961 217983 190989
rect 218011 190961 233157 190989
rect 233185 190961 233219 190989
rect 233247 190961 233281 190989
rect 233309 190961 233343 190989
rect 233371 190961 248517 190989
rect 248545 190961 248579 190989
rect 248607 190961 248641 190989
rect 248669 190961 248703 190989
rect 248731 190961 263877 190989
rect 263905 190961 263939 190989
rect 263967 190961 264001 190989
rect 264029 190961 264063 190989
rect 264091 190961 279237 190989
rect 279265 190961 279299 190989
rect 279327 190961 279361 190989
rect 279389 190961 279423 190989
rect 279451 190961 294597 190989
rect 294625 190961 294659 190989
rect 294687 190961 294721 190989
rect 294749 190961 294783 190989
rect 294811 190961 298248 190989
rect 298276 190961 298310 190989
rect 298338 190961 298372 190989
rect 298400 190961 298434 190989
rect 298462 190961 298990 190989
rect -958 190913 298990 190961
rect -958 185175 298990 185223
rect -958 185147 -910 185175
rect -882 185147 -848 185175
rect -820 185147 -786 185175
rect -758 185147 -724 185175
rect -696 185147 4617 185175
rect 4645 185147 4679 185175
rect 4707 185147 4741 185175
rect 4769 185147 4803 185175
rect 4831 185147 29939 185175
rect 29967 185147 30001 185175
rect 30029 185147 45299 185175
rect 45327 185147 45361 185175
rect 45389 185147 60659 185175
rect 60687 185147 60721 185175
rect 60749 185147 76019 185175
rect 76047 185147 76081 185175
rect 76109 185147 96777 185175
rect 96805 185147 96839 185175
rect 96867 185147 96901 185175
rect 96929 185147 96963 185175
rect 96991 185147 109939 185175
rect 109967 185147 110001 185175
rect 110029 185147 125299 185175
rect 125327 185147 125361 185175
rect 125389 185147 140659 185175
rect 140687 185147 140721 185175
rect 140749 185147 156019 185175
rect 156047 185147 156081 185175
rect 156109 185147 173577 185175
rect 173605 185147 173639 185175
rect 173667 185147 173701 185175
rect 173729 185147 173763 185175
rect 173791 185147 189939 185175
rect 189967 185147 190001 185175
rect 190029 185147 204297 185175
rect 204325 185147 204359 185175
rect 204387 185147 204421 185175
rect 204449 185147 204483 185175
rect 204511 185147 219657 185175
rect 219685 185147 219719 185175
rect 219747 185147 219781 185175
rect 219809 185147 219843 185175
rect 219871 185147 235017 185175
rect 235045 185147 235079 185175
rect 235107 185147 235141 185175
rect 235169 185147 235203 185175
rect 235231 185147 244939 185175
rect 244967 185147 245001 185175
rect 245029 185147 265737 185175
rect 265765 185147 265799 185175
rect 265827 185147 265861 185175
rect 265889 185147 265923 185175
rect 265951 185147 281097 185175
rect 281125 185147 281159 185175
rect 281187 185147 281221 185175
rect 281249 185147 281283 185175
rect 281311 185147 296457 185175
rect 296485 185147 296519 185175
rect 296547 185147 296581 185175
rect 296609 185147 296643 185175
rect 296671 185147 298728 185175
rect 298756 185147 298790 185175
rect 298818 185147 298852 185175
rect 298880 185147 298914 185175
rect 298942 185147 298990 185175
rect -958 185113 298990 185147
rect -958 185085 -910 185113
rect -882 185085 -848 185113
rect -820 185085 -786 185113
rect -758 185085 -724 185113
rect -696 185085 4617 185113
rect 4645 185085 4679 185113
rect 4707 185085 4741 185113
rect 4769 185085 4803 185113
rect 4831 185085 29939 185113
rect 29967 185085 30001 185113
rect 30029 185085 45299 185113
rect 45327 185085 45361 185113
rect 45389 185085 60659 185113
rect 60687 185085 60721 185113
rect 60749 185085 76019 185113
rect 76047 185085 76081 185113
rect 76109 185085 96777 185113
rect 96805 185085 96839 185113
rect 96867 185085 96901 185113
rect 96929 185085 96963 185113
rect 96991 185085 109939 185113
rect 109967 185085 110001 185113
rect 110029 185085 125299 185113
rect 125327 185085 125361 185113
rect 125389 185085 140659 185113
rect 140687 185085 140721 185113
rect 140749 185085 156019 185113
rect 156047 185085 156081 185113
rect 156109 185085 173577 185113
rect 173605 185085 173639 185113
rect 173667 185085 173701 185113
rect 173729 185085 173763 185113
rect 173791 185085 189939 185113
rect 189967 185085 190001 185113
rect 190029 185085 204297 185113
rect 204325 185085 204359 185113
rect 204387 185085 204421 185113
rect 204449 185085 204483 185113
rect 204511 185085 219657 185113
rect 219685 185085 219719 185113
rect 219747 185085 219781 185113
rect 219809 185085 219843 185113
rect 219871 185085 235017 185113
rect 235045 185085 235079 185113
rect 235107 185085 235141 185113
rect 235169 185085 235203 185113
rect 235231 185085 244939 185113
rect 244967 185085 245001 185113
rect 245029 185085 265737 185113
rect 265765 185085 265799 185113
rect 265827 185085 265861 185113
rect 265889 185085 265923 185113
rect 265951 185085 281097 185113
rect 281125 185085 281159 185113
rect 281187 185085 281221 185113
rect 281249 185085 281283 185113
rect 281311 185085 296457 185113
rect 296485 185085 296519 185113
rect 296547 185085 296581 185113
rect 296609 185085 296643 185113
rect 296671 185085 298728 185113
rect 298756 185085 298790 185113
rect 298818 185085 298852 185113
rect 298880 185085 298914 185113
rect 298942 185085 298990 185113
rect -958 185051 298990 185085
rect -958 185023 -910 185051
rect -882 185023 -848 185051
rect -820 185023 -786 185051
rect -758 185023 -724 185051
rect -696 185023 4617 185051
rect 4645 185023 4679 185051
rect 4707 185023 4741 185051
rect 4769 185023 4803 185051
rect 4831 185023 29939 185051
rect 29967 185023 30001 185051
rect 30029 185023 45299 185051
rect 45327 185023 45361 185051
rect 45389 185023 60659 185051
rect 60687 185023 60721 185051
rect 60749 185023 76019 185051
rect 76047 185023 76081 185051
rect 76109 185023 96777 185051
rect 96805 185023 96839 185051
rect 96867 185023 96901 185051
rect 96929 185023 96963 185051
rect 96991 185023 109939 185051
rect 109967 185023 110001 185051
rect 110029 185023 125299 185051
rect 125327 185023 125361 185051
rect 125389 185023 140659 185051
rect 140687 185023 140721 185051
rect 140749 185023 156019 185051
rect 156047 185023 156081 185051
rect 156109 185023 173577 185051
rect 173605 185023 173639 185051
rect 173667 185023 173701 185051
rect 173729 185023 173763 185051
rect 173791 185023 189939 185051
rect 189967 185023 190001 185051
rect 190029 185023 204297 185051
rect 204325 185023 204359 185051
rect 204387 185023 204421 185051
rect 204449 185023 204483 185051
rect 204511 185023 219657 185051
rect 219685 185023 219719 185051
rect 219747 185023 219781 185051
rect 219809 185023 219843 185051
rect 219871 185023 235017 185051
rect 235045 185023 235079 185051
rect 235107 185023 235141 185051
rect 235169 185023 235203 185051
rect 235231 185023 244939 185051
rect 244967 185023 245001 185051
rect 245029 185023 265737 185051
rect 265765 185023 265799 185051
rect 265827 185023 265861 185051
rect 265889 185023 265923 185051
rect 265951 185023 281097 185051
rect 281125 185023 281159 185051
rect 281187 185023 281221 185051
rect 281249 185023 281283 185051
rect 281311 185023 296457 185051
rect 296485 185023 296519 185051
rect 296547 185023 296581 185051
rect 296609 185023 296643 185051
rect 296671 185023 298728 185051
rect 298756 185023 298790 185051
rect 298818 185023 298852 185051
rect 298880 185023 298914 185051
rect 298942 185023 298990 185051
rect -958 184989 298990 185023
rect -958 184961 -910 184989
rect -882 184961 -848 184989
rect -820 184961 -786 184989
rect -758 184961 -724 184989
rect -696 184961 4617 184989
rect 4645 184961 4679 184989
rect 4707 184961 4741 184989
rect 4769 184961 4803 184989
rect 4831 184961 29939 184989
rect 29967 184961 30001 184989
rect 30029 184961 45299 184989
rect 45327 184961 45361 184989
rect 45389 184961 60659 184989
rect 60687 184961 60721 184989
rect 60749 184961 76019 184989
rect 76047 184961 76081 184989
rect 76109 184961 96777 184989
rect 96805 184961 96839 184989
rect 96867 184961 96901 184989
rect 96929 184961 96963 184989
rect 96991 184961 109939 184989
rect 109967 184961 110001 184989
rect 110029 184961 125299 184989
rect 125327 184961 125361 184989
rect 125389 184961 140659 184989
rect 140687 184961 140721 184989
rect 140749 184961 156019 184989
rect 156047 184961 156081 184989
rect 156109 184961 173577 184989
rect 173605 184961 173639 184989
rect 173667 184961 173701 184989
rect 173729 184961 173763 184989
rect 173791 184961 189939 184989
rect 189967 184961 190001 184989
rect 190029 184961 204297 184989
rect 204325 184961 204359 184989
rect 204387 184961 204421 184989
rect 204449 184961 204483 184989
rect 204511 184961 219657 184989
rect 219685 184961 219719 184989
rect 219747 184961 219781 184989
rect 219809 184961 219843 184989
rect 219871 184961 235017 184989
rect 235045 184961 235079 184989
rect 235107 184961 235141 184989
rect 235169 184961 235203 184989
rect 235231 184961 244939 184989
rect 244967 184961 245001 184989
rect 245029 184961 265737 184989
rect 265765 184961 265799 184989
rect 265827 184961 265861 184989
rect 265889 184961 265923 184989
rect 265951 184961 281097 184989
rect 281125 184961 281159 184989
rect 281187 184961 281221 184989
rect 281249 184961 281283 184989
rect 281311 184961 296457 184989
rect 296485 184961 296519 184989
rect 296547 184961 296581 184989
rect 296609 184961 296643 184989
rect 296671 184961 298728 184989
rect 298756 184961 298790 184989
rect 298818 184961 298852 184989
rect 298880 184961 298914 184989
rect 298942 184961 298990 184989
rect -958 184913 298990 184961
rect -958 182175 298990 182223
rect -958 182147 -430 182175
rect -402 182147 -368 182175
rect -340 182147 -306 182175
rect -278 182147 -244 182175
rect -216 182147 2757 182175
rect 2785 182147 2819 182175
rect 2847 182147 2881 182175
rect 2909 182147 2943 182175
rect 2971 182147 18117 182175
rect 18145 182147 18179 182175
rect 18207 182147 18241 182175
rect 18269 182147 18303 182175
rect 18331 182147 22259 182175
rect 22287 182147 22321 182175
rect 22349 182147 37619 182175
rect 37647 182147 37681 182175
rect 37709 182147 52979 182175
rect 53007 182147 53041 182175
rect 53069 182147 68339 182175
rect 68367 182147 68401 182175
rect 68429 182147 83699 182175
rect 83727 182147 83761 182175
rect 83789 182147 94917 182175
rect 94945 182147 94979 182175
rect 95007 182147 95041 182175
rect 95069 182147 95103 182175
rect 95131 182147 102259 182175
rect 102287 182147 102321 182175
rect 102349 182147 117619 182175
rect 117647 182147 117681 182175
rect 117709 182147 132979 182175
rect 133007 182147 133041 182175
rect 133069 182147 148339 182175
rect 148367 182147 148401 182175
rect 148429 182147 163699 182175
rect 163727 182147 163761 182175
rect 163789 182147 171717 182175
rect 171745 182147 171779 182175
rect 171807 182147 171841 182175
rect 171869 182147 171903 182175
rect 171931 182147 182259 182175
rect 182287 182147 182321 182175
rect 182349 182147 197619 182175
rect 197647 182147 197681 182175
rect 197709 182147 202437 182175
rect 202465 182147 202499 182175
rect 202527 182147 202561 182175
rect 202589 182147 202623 182175
rect 202651 182147 217797 182175
rect 217825 182147 217859 182175
rect 217887 182147 217921 182175
rect 217949 182147 217983 182175
rect 218011 182147 233157 182175
rect 233185 182147 233219 182175
rect 233247 182147 233281 182175
rect 233309 182147 233343 182175
rect 233371 182147 237259 182175
rect 237287 182147 237321 182175
rect 237349 182147 252619 182175
rect 252647 182147 252681 182175
rect 252709 182147 263877 182175
rect 263905 182147 263939 182175
rect 263967 182147 264001 182175
rect 264029 182147 264063 182175
rect 264091 182147 279237 182175
rect 279265 182147 279299 182175
rect 279327 182147 279361 182175
rect 279389 182147 279423 182175
rect 279451 182147 294597 182175
rect 294625 182147 294659 182175
rect 294687 182147 294721 182175
rect 294749 182147 294783 182175
rect 294811 182147 298248 182175
rect 298276 182147 298310 182175
rect 298338 182147 298372 182175
rect 298400 182147 298434 182175
rect 298462 182147 298990 182175
rect -958 182113 298990 182147
rect -958 182085 -430 182113
rect -402 182085 -368 182113
rect -340 182085 -306 182113
rect -278 182085 -244 182113
rect -216 182085 2757 182113
rect 2785 182085 2819 182113
rect 2847 182085 2881 182113
rect 2909 182085 2943 182113
rect 2971 182085 18117 182113
rect 18145 182085 18179 182113
rect 18207 182085 18241 182113
rect 18269 182085 18303 182113
rect 18331 182085 22259 182113
rect 22287 182085 22321 182113
rect 22349 182085 37619 182113
rect 37647 182085 37681 182113
rect 37709 182085 52979 182113
rect 53007 182085 53041 182113
rect 53069 182085 68339 182113
rect 68367 182085 68401 182113
rect 68429 182085 83699 182113
rect 83727 182085 83761 182113
rect 83789 182085 94917 182113
rect 94945 182085 94979 182113
rect 95007 182085 95041 182113
rect 95069 182085 95103 182113
rect 95131 182085 102259 182113
rect 102287 182085 102321 182113
rect 102349 182085 117619 182113
rect 117647 182085 117681 182113
rect 117709 182085 132979 182113
rect 133007 182085 133041 182113
rect 133069 182085 148339 182113
rect 148367 182085 148401 182113
rect 148429 182085 163699 182113
rect 163727 182085 163761 182113
rect 163789 182085 171717 182113
rect 171745 182085 171779 182113
rect 171807 182085 171841 182113
rect 171869 182085 171903 182113
rect 171931 182085 182259 182113
rect 182287 182085 182321 182113
rect 182349 182085 197619 182113
rect 197647 182085 197681 182113
rect 197709 182085 202437 182113
rect 202465 182085 202499 182113
rect 202527 182085 202561 182113
rect 202589 182085 202623 182113
rect 202651 182085 217797 182113
rect 217825 182085 217859 182113
rect 217887 182085 217921 182113
rect 217949 182085 217983 182113
rect 218011 182085 233157 182113
rect 233185 182085 233219 182113
rect 233247 182085 233281 182113
rect 233309 182085 233343 182113
rect 233371 182085 237259 182113
rect 237287 182085 237321 182113
rect 237349 182085 252619 182113
rect 252647 182085 252681 182113
rect 252709 182085 263877 182113
rect 263905 182085 263939 182113
rect 263967 182085 264001 182113
rect 264029 182085 264063 182113
rect 264091 182085 279237 182113
rect 279265 182085 279299 182113
rect 279327 182085 279361 182113
rect 279389 182085 279423 182113
rect 279451 182085 294597 182113
rect 294625 182085 294659 182113
rect 294687 182085 294721 182113
rect 294749 182085 294783 182113
rect 294811 182085 298248 182113
rect 298276 182085 298310 182113
rect 298338 182085 298372 182113
rect 298400 182085 298434 182113
rect 298462 182085 298990 182113
rect -958 182051 298990 182085
rect -958 182023 -430 182051
rect -402 182023 -368 182051
rect -340 182023 -306 182051
rect -278 182023 -244 182051
rect -216 182023 2757 182051
rect 2785 182023 2819 182051
rect 2847 182023 2881 182051
rect 2909 182023 2943 182051
rect 2971 182023 18117 182051
rect 18145 182023 18179 182051
rect 18207 182023 18241 182051
rect 18269 182023 18303 182051
rect 18331 182023 22259 182051
rect 22287 182023 22321 182051
rect 22349 182023 37619 182051
rect 37647 182023 37681 182051
rect 37709 182023 52979 182051
rect 53007 182023 53041 182051
rect 53069 182023 68339 182051
rect 68367 182023 68401 182051
rect 68429 182023 83699 182051
rect 83727 182023 83761 182051
rect 83789 182023 94917 182051
rect 94945 182023 94979 182051
rect 95007 182023 95041 182051
rect 95069 182023 95103 182051
rect 95131 182023 102259 182051
rect 102287 182023 102321 182051
rect 102349 182023 117619 182051
rect 117647 182023 117681 182051
rect 117709 182023 132979 182051
rect 133007 182023 133041 182051
rect 133069 182023 148339 182051
rect 148367 182023 148401 182051
rect 148429 182023 163699 182051
rect 163727 182023 163761 182051
rect 163789 182023 171717 182051
rect 171745 182023 171779 182051
rect 171807 182023 171841 182051
rect 171869 182023 171903 182051
rect 171931 182023 182259 182051
rect 182287 182023 182321 182051
rect 182349 182023 197619 182051
rect 197647 182023 197681 182051
rect 197709 182023 202437 182051
rect 202465 182023 202499 182051
rect 202527 182023 202561 182051
rect 202589 182023 202623 182051
rect 202651 182023 217797 182051
rect 217825 182023 217859 182051
rect 217887 182023 217921 182051
rect 217949 182023 217983 182051
rect 218011 182023 233157 182051
rect 233185 182023 233219 182051
rect 233247 182023 233281 182051
rect 233309 182023 233343 182051
rect 233371 182023 237259 182051
rect 237287 182023 237321 182051
rect 237349 182023 252619 182051
rect 252647 182023 252681 182051
rect 252709 182023 263877 182051
rect 263905 182023 263939 182051
rect 263967 182023 264001 182051
rect 264029 182023 264063 182051
rect 264091 182023 279237 182051
rect 279265 182023 279299 182051
rect 279327 182023 279361 182051
rect 279389 182023 279423 182051
rect 279451 182023 294597 182051
rect 294625 182023 294659 182051
rect 294687 182023 294721 182051
rect 294749 182023 294783 182051
rect 294811 182023 298248 182051
rect 298276 182023 298310 182051
rect 298338 182023 298372 182051
rect 298400 182023 298434 182051
rect 298462 182023 298990 182051
rect -958 181989 298990 182023
rect -958 181961 -430 181989
rect -402 181961 -368 181989
rect -340 181961 -306 181989
rect -278 181961 -244 181989
rect -216 181961 2757 181989
rect 2785 181961 2819 181989
rect 2847 181961 2881 181989
rect 2909 181961 2943 181989
rect 2971 181961 18117 181989
rect 18145 181961 18179 181989
rect 18207 181961 18241 181989
rect 18269 181961 18303 181989
rect 18331 181961 22259 181989
rect 22287 181961 22321 181989
rect 22349 181961 37619 181989
rect 37647 181961 37681 181989
rect 37709 181961 52979 181989
rect 53007 181961 53041 181989
rect 53069 181961 68339 181989
rect 68367 181961 68401 181989
rect 68429 181961 83699 181989
rect 83727 181961 83761 181989
rect 83789 181961 94917 181989
rect 94945 181961 94979 181989
rect 95007 181961 95041 181989
rect 95069 181961 95103 181989
rect 95131 181961 102259 181989
rect 102287 181961 102321 181989
rect 102349 181961 117619 181989
rect 117647 181961 117681 181989
rect 117709 181961 132979 181989
rect 133007 181961 133041 181989
rect 133069 181961 148339 181989
rect 148367 181961 148401 181989
rect 148429 181961 163699 181989
rect 163727 181961 163761 181989
rect 163789 181961 171717 181989
rect 171745 181961 171779 181989
rect 171807 181961 171841 181989
rect 171869 181961 171903 181989
rect 171931 181961 182259 181989
rect 182287 181961 182321 181989
rect 182349 181961 197619 181989
rect 197647 181961 197681 181989
rect 197709 181961 202437 181989
rect 202465 181961 202499 181989
rect 202527 181961 202561 181989
rect 202589 181961 202623 181989
rect 202651 181961 217797 181989
rect 217825 181961 217859 181989
rect 217887 181961 217921 181989
rect 217949 181961 217983 181989
rect 218011 181961 233157 181989
rect 233185 181961 233219 181989
rect 233247 181961 233281 181989
rect 233309 181961 233343 181989
rect 233371 181961 237259 181989
rect 237287 181961 237321 181989
rect 237349 181961 252619 181989
rect 252647 181961 252681 181989
rect 252709 181961 263877 181989
rect 263905 181961 263939 181989
rect 263967 181961 264001 181989
rect 264029 181961 264063 181989
rect 264091 181961 279237 181989
rect 279265 181961 279299 181989
rect 279327 181961 279361 181989
rect 279389 181961 279423 181989
rect 279451 181961 294597 181989
rect 294625 181961 294659 181989
rect 294687 181961 294721 181989
rect 294749 181961 294783 181989
rect 294811 181961 298248 181989
rect 298276 181961 298310 181989
rect 298338 181961 298372 181989
rect 298400 181961 298434 181989
rect 298462 181961 298990 181989
rect -958 181913 298990 181961
rect -958 176175 298990 176223
rect -958 176147 -910 176175
rect -882 176147 -848 176175
rect -820 176147 -786 176175
rect -758 176147 -724 176175
rect -696 176147 4617 176175
rect 4645 176147 4679 176175
rect 4707 176147 4741 176175
rect 4769 176147 4803 176175
rect 4831 176147 29939 176175
rect 29967 176147 30001 176175
rect 30029 176147 45299 176175
rect 45327 176147 45361 176175
rect 45389 176147 60659 176175
rect 60687 176147 60721 176175
rect 60749 176147 76019 176175
rect 76047 176147 76081 176175
rect 76109 176147 96777 176175
rect 96805 176147 96839 176175
rect 96867 176147 96901 176175
rect 96929 176147 96963 176175
rect 96991 176147 109939 176175
rect 109967 176147 110001 176175
rect 110029 176147 125299 176175
rect 125327 176147 125361 176175
rect 125389 176147 140659 176175
rect 140687 176147 140721 176175
rect 140749 176147 156019 176175
rect 156047 176147 156081 176175
rect 156109 176147 173577 176175
rect 173605 176147 173639 176175
rect 173667 176147 173701 176175
rect 173729 176147 173763 176175
rect 173791 176147 189939 176175
rect 189967 176147 190001 176175
rect 190029 176147 204297 176175
rect 204325 176147 204359 176175
rect 204387 176147 204421 176175
rect 204449 176147 204483 176175
rect 204511 176147 219657 176175
rect 219685 176147 219719 176175
rect 219747 176147 219781 176175
rect 219809 176147 219843 176175
rect 219871 176147 235017 176175
rect 235045 176147 235079 176175
rect 235107 176147 235141 176175
rect 235169 176147 235203 176175
rect 235231 176147 244939 176175
rect 244967 176147 245001 176175
rect 245029 176147 265737 176175
rect 265765 176147 265799 176175
rect 265827 176147 265861 176175
rect 265889 176147 265923 176175
rect 265951 176147 281097 176175
rect 281125 176147 281159 176175
rect 281187 176147 281221 176175
rect 281249 176147 281283 176175
rect 281311 176147 296457 176175
rect 296485 176147 296519 176175
rect 296547 176147 296581 176175
rect 296609 176147 296643 176175
rect 296671 176147 298728 176175
rect 298756 176147 298790 176175
rect 298818 176147 298852 176175
rect 298880 176147 298914 176175
rect 298942 176147 298990 176175
rect -958 176113 298990 176147
rect -958 176085 -910 176113
rect -882 176085 -848 176113
rect -820 176085 -786 176113
rect -758 176085 -724 176113
rect -696 176085 4617 176113
rect 4645 176085 4679 176113
rect 4707 176085 4741 176113
rect 4769 176085 4803 176113
rect 4831 176085 29939 176113
rect 29967 176085 30001 176113
rect 30029 176085 45299 176113
rect 45327 176085 45361 176113
rect 45389 176085 60659 176113
rect 60687 176085 60721 176113
rect 60749 176085 76019 176113
rect 76047 176085 76081 176113
rect 76109 176085 96777 176113
rect 96805 176085 96839 176113
rect 96867 176085 96901 176113
rect 96929 176085 96963 176113
rect 96991 176085 109939 176113
rect 109967 176085 110001 176113
rect 110029 176085 125299 176113
rect 125327 176085 125361 176113
rect 125389 176085 140659 176113
rect 140687 176085 140721 176113
rect 140749 176085 156019 176113
rect 156047 176085 156081 176113
rect 156109 176085 173577 176113
rect 173605 176085 173639 176113
rect 173667 176085 173701 176113
rect 173729 176085 173763 176113
rect 173791 176085 189939 176113
rect 189967 176085 190001 176113
rect 190029 176085 204297 176113
rect 204325 176085 204359 176113
rect 204387 176085 204421 176113
rect 204449 176085 204483 176113
rect 204511 176085 219657 176113
rect 219685 176085 219719 176113
rect 219747 176085 219781 176113
rect 219809 176085 219843 176113
rect 219871 176085 235017 176113
rect 235045 176085 235079 176113
rect 235107 176085 235141 176113
rect 235169 176085 235203 176113
rect 235231 176085 244939 176113
rect 244967 176085 245001 176113
rect 245029 176085 265737 176113
rect 265765 176085 265799 176113
rect 265827 176085 265861 176113
rect 265889 176085 265923 176113
rect 265951 176085 281097 176113
rect 281125 176085 281159 176113
rect 281187 176085 281221 176113
rect 281249 176085 281283 176113
rect 281311 176085 296457 176113
rect 296485 176085 296519 176113
rect 296547 176085 296581 176113
rect 296609 176085 296643 176113
rect 296671 176085 298728 176113
rect 298756 176085 298790 176113
rect 298818 176085 298852 176113
rect 298880 176085 298914 176113
rect 298942 176085 298990 176113
rect -958 176051 298990 176085
rect -958 176023 -910 176051
rect -882 176023 -848 176051
rect -820 176023 -786 176051
rect -758 176023 -724 176051
rect -696 176023 4617 176051
rect 4645 176023 4679 176051
rect 4707 176023 4741 176051
rect 4769 176023 4803 176051
rect 4831 176023 29939 176051
rect 29967 176023 30001 176051
rect 30029 176023 45299 176051
rect 45327 176023 45361 176051
rect 45389 176023 60659 176051
rect 60687 176023 60721 176051
rect 60749 176023 76019 176051
rect 76047 176023 76081 176051
rect 76109 176023 96777 176051
rect 96805 176023 96839 176051
rect 96867 176023 96901 176051
rect 96929 176023 96963 176051
rect 96991 176023 109939 176051
rect 109967 176023 110001 176051
rect 110029 176023 125299 176051
rect 125327 176023 125361 176051
rect 125389 176023 140659 176051
rect 140687 176023 140721 176051
rect 140749 176023 156019 176051
rect 156047 176023 156081 176051
rect 156109 176023 173577 176051
rect 173605 176023 173639 176051
rect 173667 176023 173701 176051
rect 173729 176023 173763 176051
rect 173791 176023 189939 176051
rect 189967 176023 190001 176051
rect 190029 176023 204297 176051
rect 204325 176023 204359 176051
rect 204387 176023 204421 176051
rect 204449 176023 204483 176051
rect 204511 176023 219657 176051
rect 219685 176023 219719 176051
rect 219747 176023 219781 176051
rect 219809 176023 219843 176051
rect 219871 176023 235017 176051
rect 235045 176023 235079 176051
rect 235107 176023 235141 176051
rect 235169 176023 235203 176051
rect 235231 176023 244939 176051
rect 244967 176023 245001 176051
rect 245029 176023 265737 176051
rect 265765 176023 265799 176051
rect 265827 176023 265861 176051
rect 265889 176023 265923 176051
rect 265951 176023 281097 176051
rect 281125 176023 281159 176051
rect 281187 176023 281221 176051
rect 281249 176023 281283 176051
rect 281311 176023 296457 176051
rect 296485 176023 296519 176051
rect 296547 176023 296581 176051
rect 296609 176023 296643 176051
rect 296671 176023 298728 176051
rect 298756 176023 298790 176051
rect 298818 176023 298852 176051
rect 298880 176023 298914 176051
rect 298942 176023 298990 176051
rect -958 175989 298990 176023
rect -958 175961 -910 175989
rect -882 175961 -848 175989
rect -820 175961 -786 175989
rect -758 175961 -724 175989
rect -696 175961 4617 175989
rect 4645 175961 4679 175989
rect 4707 175961 4741 175989
rect 4769 175961 4803 175989
rect 4831 175961 29939 175989
rect 29967 175961 30001 175989
rect 30029 175961 45299 175989
rect 45327 175961 45361 175989
rect 45389 175961 60659 175989
rect 60687 175961 60721 175989
rect 60749 175961 76019 175989
rect 76047 175961 76081 175989
rect 76109 175961 96777 175989
rect 96805 175961 96839 175989
rect 96867 175961 96901 175989
rect 96929 175961 96963 175989
rect 96991 175961 109939 175989
rect 109967 175961 110001 175989
rect 110029 175961 125299 175989
rect 125327 175961 125361 175989
rect 125389 175961 140659 175989
rect 140687 175961 140721 175989
rect 140749 175961 156019 175989
rect 156047 175961 156081 175989
rect 156109 175961 173577 175989
rect 173605 175961 173639 175989
rect 173667 175961 173701 175989
rect 173729 175961 173763 175989
rect 173791 175961 189939 175989
rect 189967 175961 190001 175989
rect 190029 175961 204297 175989
rect 204325 175961 204359 175989
rect 204387 175961 204421 175989
rect 204449 175961 204483 175989
rect 204511 175961 219657 175989
rect 219685 175961 219719 175989
rect 219747 175961 219781 175989
rect 219809 175961 219843 175989
rect 219871 175961 235017 175989
rect 235045 175961 235079 175989
rect 235107 175961 235141 175989
rect 235169 175961 235203 175989
rect 235231 175961 244939 175989
rect 244967 175961 245001 175989
rect 245029 175961 265737 175989
rect 265765 175961 265799 175989
rect 265827 175961 265861 175989
rect 265889 175961 265923 175989
rect 265951 175961 281097 175989
rect 281125 175961 281159 175989
rect 281187 175961 281221 175989
rect 281249 175961 281283 175989
rect 281311 175961 296457 175989
rect 296485 175961 296519 175989
rect 296547 175961 296581 175989
rect 296609 175961 296643 175989
rect 296671 175961 298728 175989
rect 298756 175961 298790 175989
rect 298818 175961 298852 175989
rect 298880 175961 298914 175989
rect 298942 175961 298990 175989
rect -958 175913 298990 175961
rect -958 173175 298990 173223
rect -958 173147 -430 173175
rect -402 173147 -368 173175
rect -340 173147 -306 173175
rect -278 173147 -244 173175
rect -216 173147 2757 173175
rect 2785 173147 2819 173175
rect 2847 173147 2881 173175
rect 2909 173147 2943 173175
rect 2971 173147 18117 173175
rect 18145 173147 18179 173175
rect 18207 173147 18241 173175
rect 18269 173147 18303 173175
rect 18331 173147 22259 173175
rect 22287 173147 22321 173175
rect 22349 173147 37619 173175
rect 37647 173147 37681 173175
rect 37709 173147 52979 173175
rect 53007 173147 53041 173175
rect 53069 173147 68339 173175
rect 68367 173147 68401 173175
rect 68429 173147 83699 173175
rect 83727 173147 83761 173175
rect 83789 173147 94917 173175
rect 94945 173147 94979 173175
rect 95007 173147 95041 173175
rect 95069 173147 95103 173175
rect 95131 173147 102259 173175
rect 102287 173147 102321 173175
rect 102349 173147 117619 173175
rect 117647 173147 117681 173175
rect 117709 173147 132979 173175
rect 133007 173147 133041 173175
rect 133069 173147 148339 173175
rect 148367 173147 148401 173175
rect 148429 173147 163699 173175
rect 163727 173147 163761 173175
rect 163789 173147 171717 173175
rect 171745 173147 171779 173175
rect 171807 173147 171841 173175
rect 171869 173147 171903 173175
rect 171931 173147 182259 173175
rect 182287 173147 182321 173175
rect 182349 173147 187077 173175
rect 187105 173147 187139 173175
rect 187167 173147 187201 173175
rect 187229 173147 187263 173175
rect 187291 173147 197619 173175
rect 197647 173147 197681 173175
rect 197709 173147 202437 173175
rect 202465 173147 202499 173175
rect 202527 173147 202561 173175
rect 202589 173147 202623 173175
rect 202651 173147 217797 173175
rect 217825 173147 217859 173175
rect 217887 173147 217921 173175
rect 217949 173147 217983 173175
rect 218011 173147 233157 173175
rect 233185 173147 233219 173175
rect 233247 173147 233281 173175
rect 233309 173147 233343 173175
rect 233371 173147 237259 173175
rect 237287 173147 237321 173175
rect 237349 173147 252619 173175
rect 252647 173147 252681 173175
rect 252709 173147 263877 173175
rect 263905 173147 263939 173175
rect 263967 173147 264001 173175
rect 264029 173147 264063 173175
rect 264091 173147 279237 173175
rect 279265 173147 279299 173175
rect 279327 173147 279361 173175
rect 279389 173147 279423 173175
rect 279451 173147 294597 173175
rect 294625 173147 294659 173175
rect 294687 173147 294721 173175
rect 294749 173147 294783 173175
rect 294811 173147 298248 173175
rect 298276 173147 298310 173175
rect 298338 173147 298372 173175
rect 298400 173147 298434 173175
rect 298462 173147 298990 173175
rect -958 173113 298990 173147
rect -958 173085 -430 173113
rect -402 173085 -368 173113
rect -340 173085 -306 173113
rect -278 173085 -244 173113
rect -216 173085 2757 173113
rect 2785 173085 2819 173113
rect 2847 173085 2881 173113
rect 2909 173085 2943 173113
rect 2971 173085 18117 173113
rect 18145 173085 18179 173113
rect 18207 173085 18241 173113
rect 18269 173085 18303 173113
rect 18331 173085 22259 173113
rect 22287 173085 22321 173113
rect 22349 173085 37619 173113
rect 37647 173085 37681 173113
rect 37709 173085 52979 173113
rect 53007 173085 53041 173113
rect 53069 173085 68339 173113
rect 68367 173085 68401 173113
rect 68429 173085 83699 173113
rect 83727 173085 83761 173113
rect 83789 173085 94917 173113
rect 94945 173085 94979 173113
rect 95007 173085 95041 173113
rect 95069 173085 95103 173113
rect 95131 173085 102259 173113
rect 102287 173085 102321 173113
rect 102349 173085 117619 173113
rect 117647 173085 117681 173113
rect 117709 173085 132979 173113
rect 133007 173085 133041 173113
rect 133069 173085 148339 173113
rect 148367 173085 148401 173113
rect 148429 173085 163699 173113
rect 163727 173085 163761 173113
rect 163789 173085 171717 173113
rect 171745 173085 171779 173113
rect 171807 173085 171841 173113
rect 171869 173085 171903 173113
rect 171931 173085 182259 173113
rect 182287 173085 182321 173113
rect 182349 173085 187077 173113
rect 187105 173085 187139 173113
rect 187167 173085 187201 173113
rect 187229 173085 187263 173113
rect 187291 173085 197619 173113
rect 197647 173085 197681 173113
rect 197709 173085 202437 173113
rect 202465 173085 202499 173113
rect 202527 173085 202561 173113
rect 202589 173085 202623 173113
rect 202651 173085 217797 173113
rect 217825 173085 217859 173113
rect 217887 173085 217921 173113
rect 217949 173085 217983 173113
rect 218011 173085 233157 173113
rect 233185 173085 233219 173113
rect 233247 173085 233281 173113
rect 233309 173085 233343 173113
rect 233371 173085 237259 173113
rect 237287 173085 237321 173113
rect 237349 173085 252619 173113
rect 252647 173085 252681 173113
rect 252709 173085 263877 173113
rect 263905 173085 263939 173113
rect 263967 173085 264001 173113
rect 264029 173085 264063 173113
rect 264091 173085 279237 173113
rect 279265 173085 279299 173113
rect 279327 173085 279361 173113
rect 279389 173085 279423 173113
rect 279451 173085 294597 173113
rect 294625 173085 294659 173113
rect 294687 173085 294721 173113
rect 294749 173085 294783 173113
rect 294811 173085 298248 173113
rect 298276 173085 298310 173113
rect 298338 173085 298372 173113
rect 298400 173085 298434 173113
rect 298462 173085 298990 173113
rect -958 173051 298990 173085
rect -958 173023 -430 173051
rect -402 173023 -368 173051
rect -340 173023 -306 173051
rect -278 173023 -244 173051
rect -216 173023 2757 173051
rect 2785 173023 2819 173051
rect 2847 173023 2881 173051
rect 2909 173023 2943 173051
rect 2971 173023 18117 173051
rect 18145 173023 18179 173051
rect 18207 173023 18241 173051
rect 18269 173023 18303 173051
rect 18331 173023 22259 173051
rect 22287 173023 22321 173051
rect 22349 173023 37619 173051
rect 37647 173023 37681 173051
rect 37709 173023 52979 173051
rect 53007 173023 53041 173051
rect 53069 173023 68339 173051
rect 68367 173023 68401 173051
rect 68429 173023 83699 173051
rect 83727 173023 83761 173051
rect 83789 173023 94917 173051
rect 94945 173023 94979 173051
rect 95007 173023 95041 173051
rect 95069 173023 95103 173051
rect 95131 173023 102259 173051
rect 102287 173023 102321 173051
rect 102349 173023 117619 173051
rect 117647 173023 117681 173051
rect 117709 173023 132979 173051
rect 133007 173023 133041 173051
rect 133069 173023 148339 173051
rect 148367 173023 148401 173051
rect 148429 173023 163699 173051
rect 163727 173023 163761 173051
rect 163789 173023 171717 173051
rect 171745 173023 171779 173051
rect 171807 173023 171841 173051
rect 171869 173023 171903 173051
rect 171931 173023 182259 173051
rect 182287 173023 182321 173051
rect 182349 173023 187077 173051
rect 187105 173023 187139 173051
rect 187167 173023 187201 173051
rect 187229 173023 187263 173051
rect 187291 173023 197619 173051
rect 197647 173023 197681 173051
rect 197709 173023 202437 173051
rect 202465 173023 202499 173051
rect 202527 173023 202561 173051
rect 202589 173023 202623 173051
rect 202651 173023 217797 173051
rect 217825 173023 217859 173051
rect 217887 173023 217921 173051
rect 217949 173023 217983 173051
rect 218011 173023 233157 173051
rect 233185 173023 233219 173051
rect 233247 173023 233281 173051
rect 233309 173023 233343 173051
rect 233371 173023 237259 173051
rect 237287 173023 237321 173051
rect 237349 173023 252619 173051
rect 252647 173023 252681 173051
rect 252709 173023 263877 173051
rect 263905 173023 263939 173051
rect 263967 173023 264001 173051
rect 264029 173023 264063 173051
rect 264091 173023 279237 173051
rect 279265 173023 279299 173051
rect 279327 173023 279361 173051
rect 279389 173023 279423 173051
rect 279451 173023 294597 173051
rect 294625 173023 294659 173051
rect 294687 173023 294721 173051
rect 294749 173023 294783 173051
rect 294811 173023 298248 173051
rect 298276 173023 298310 173051
rect 298338 173023 298372 173051
rect 298400 173023 298434 173051
rect 298462 173023 298990 173051
rect -958 172989 298990 173023
rect -958 172961 -430 172989
rect -402 172961 -368 172989
rect -340 172961 -306 172989
rect -278 172961 -244 172989
rect -216 172961 2757 172989
rect 2785 172961 2819 172989
rect 2847 172961 2881 172989
rect 2909 172961 2943 172989
rect 2971 172961 18117 172989
rect 18145 172961 18179 172989
rect 18207 172961 18241 172989
rect 18269 172961 18303 172989
rect 18331 172961 22259 172989
rect 22287 172961 22321 172989
rect 22349 172961 37619 172989
rect 37647 172961 37681 172989
rect 37709 172961 52979 172989
rect 53007 172961 53041 172989
rect 53069 172961 68339 172989
rect 68367 172961 68401 172989
rect 68429 172961 83699 172989
rect 83727 172961 83761 172989
rect 83789 172961 94917 172989
rect 94945 172961 94979 172989
rect 95007 172961 95041 172989
rect 95069 172961 95103 172989
rect 95131 172961 102259 172989
rect 102287 172961 102321 172989
rect 102349 172961 117619 172989
rect 117647 172961 117681 172989
rect 117709 172961 132979 172989
rect 133007 172961 133041 172989
rect 133069 172961 148339 172989
rect 148367 172961 148401 172989
rect 148429 172961 163699 172989
rect 163727 172961 163761 172989
rect 163789 172961 171717 172989
rect 171745 172961 171779 172989
rect 171807 172961 171841 172989
rect 171869 172961 171903 172989
rect 171931 172961 182259 172989
rect 182287 172961 182321 172989
rect 182349 172961 187077 172989
rect 187105 172961 187139 172989
rect 187167 172961 187201 172989
rect 187229 172961 187263 172989
rect 187291 172961 197619 172989
rect 197647 172961 197681 172989
rect 197709 172961 202437 172989
rect 202465 172961 202499 172989
rect 202527 172961 202561 172989
rect 202589 172961 202623 172989
rect 202651 172961 217797 172989
rect 217825 172961 217859 172989
rect 217887 172961 217921 172989
rect 217949 172961 217983 172989
rect 218011 172961 233157 172989
rect 233185 172961 233219 172989
rect 233247 172961 233281 172989
rect 233309 172961 233343 172989
rect 233371 172961 237259 172989
rect 237287 172961 237321 172989
rect 237349 172961 252619 172989
rect 252647 172961 252681 172989
rect 252709 172961 263877 172989
rect 263905 172961 263939 172989
rect 263967 172961 264001 172989
rect 264029 172961 264063 172989
rect 264091 172961 279237 172989
rect 279265 172961 279299 172989
rect 279327 172961 279361 172989
rect 279389 172961 279423 172989
rect 279451 172961 294597 172989
rect 294625 172961 294659 172989
rect 294687 172961 294721 172989
rect 294749 172961 294783 172989
rect 294811 172961 298248 172989
rect 298276 172961 298310 172989
rect 298338 172961 298372 172989
rect 298400 172961 298434 172989
rect 298462 172961 298990 172989
rect -958 172913 298990 172961
rect -958 167175 298990 167223
rect -958 167147 -910 167175
rect -882 167147 -848 167175
rect -820 167147 -786 167175
rect -758 167147 -724 167175
rect -696 167147 4617 167175
rect 4645 167147 4679 167175
rect 4707 167147 4741 167175
rect 4769 167147 4803 167175
rect 4831 167147 19977 167175
rect 20005 167147 20039 167175
rect 20067 167147 20101 167175
rect 20129 167147 20163 167175
rect 20191 167147 35337 167175
rect 35365 167147 35399 167175
rect 35427 167147 35461 167175
rect 35489 167147 35523 167175
rect 35551 167147 50697 167175
rect 50725 167147 50759 167175
rect 50787 167147 50821 167175
rect 50849 167147 50883 167175
rect 50911 167147 66057 167175
rect 66085 167147 66119 167175
rect 66147 167147 66181 167175
rect 66209 167147 66243 167175
rect 66271 167147 81417 167175
rect 81445 167147 81479 167175
rect 81507 167147 81541 167175
rect 81569 167147 81603 167175
rect 81631 167147 96777 167175
rect 96805 167147 96839 167175
rect 96867 167147 96901 167175
rect 96929 167147 96963 167175
rect 96991 167147 173577 167175
rect 173605 167147 173639 167175
rect 173667 167147 173701 167175
rect 173729 167147 173763 167175
rect 173791 167147 204297 167175
rect 204325 167147 204359 167175
rect 204387 167147 204421 167175
rect 204449 167147 204483 167175
rect 204511 167147 219657 167175
rect 219685 167147 219719 167175
rect 219747 167147 219781 167175
rect 219809 167147 219843 167175
rect 219871 167147 235017 167175
rect 235045 167147 235079 167175
rect 235107 167147 235141 167175
rect 235169 167147 235203 167175
rect 235231 167147 250377 167175
rect 250405 167147 250439 167175
rect 250467 167147 250501 167175
rect 250529 167147 250563 167175
rect 250591 167147 265737 167175
rect 265765 167147 265799 167175
rect 265827 167147 265861 167175
rect 265889 167147 265923 167175
rect 265951 167147 281097 167175
rect 281125 167147 281159 167175
rect 281187 167147 281221 167175
rect 281249 167147 281283 167175
rect 281311 167147 296457 167175
rect 296485 167147 296519 167175
rect 296547 167147 296581 167175
rect 296609 167147 296643 167175
rect 296671 167147 298728 167175
rect 298756 167147 298790 167175
rect 298818 167147 298852 167175
rect 298880 167147 298914 167175
rect 298942 167147 298990 167175
rect -958 167113 298990 167147
rect -958 167085 -910 167113
rect -882 167085 -848 167113
rect -820 167085 -786 167113
rect -758 167085 -724 167113
rect -696 167085 4617 167113
rect 4645 167085 4679 167113
rect 4707 167085 4741 167113
rect 4769 167085 4803 167113
rect 4831 167085 19977 167113
rect 20005 167085 20039 167113
rect 20067 167085 20101 167113
rect 20129 167085 20163 167113
rect 20191 167085 35337 167113
rect 35365 167085 35399 167113
rect 35427 167085 35461 167113
rect 35489 167085 35523 167113
rect 35551 167085 50697 167113
rect 50725 167085 50759 167113
rect 50787 167085 50821 167113
rect 50849 167085 50883 167113
rect 50911 167085 66057 167113
rect 66085 167085 66119 167113
rect 66147 167085 66181 167113
rect 66209 167085 66243 167113
rect 66271 167085 81417 167113
rect 81445 167085 81479 167113
rect 81507 167085 81541 167113
rect 81569 167085 81603 167113
rect 81631 167085 96777 167113
rect 96805 167085 96839 167113
rect 96867 167085 96901 167113
rect 96929 167085 96963 167113
rect 96991 167085 173577 167113
rect 173605 167085 173639 167113
rect 173667 167085 173701 167113
rect 173729 167085 173763 167113
rect 173791 167085 204297 167113
rect 204325 167085 204359 167113
rect 204387 167085 204421 167113
rect 204449 167085 204483 167113
rect 204511 167085 219657 167113
rect 219685 167085 219719 167113
rect 219747 167085 219781 167113
rect 219809 167085 219843 167113
rect 219871 167085 235017 167113
rect 235045 167085 235079 167113
rect 235107 167085 235141 167113
rect 235169 167085 235203 167113
rect 235231 167085 250377 167113
rect 250405 167085 250439 167113
rect 250467 167085 250501 167113
rect 250529 167085 250563 167113
rect 250591 167085 265737 167113
rect 265765 167085 265799 167113
rect 265827 167085 265861 167113
rect 265889 167085 265923 167113
rect 265951 167085 281097 167113
rect 281125 167085 281159 167113
rect 281187 167085 281221 167113
rect 281249 167085 281283 167113
rect 281311 167085 296457 167113
rect 296485 167085 296519 167113
rect 296547 167085 296581 167113
rect 296609 167085 296643 167113
rect 296671 167085 298728 167113
rect 298756 167085 298790 167113
rect 298818 167085 298852 167113
rect 298880 167085 298914 167113
rect 298942 167085 298990 167113
rect -958 167051 298990 167085
rect -958 167023 -910 167051
rect -882 167023 -848 167051
rect -820 167023 -786 167051
rect -758 167023 -724 167051
rect -696 167023 4617 167051
rect 4645 167023 4679 167051
rect 4707 167023 4741 167051
rect 4769 167023 4803 167051
rect 4831 167023 19977 167051
rect 20005 167023 20039 167051
rect 20067 167023 20101 167051
rect 20129 167023 20163 167051
rect 20191 167023 35337 167051
rect 35365 167023 35399 167051
rect 35427 167023 35461 167051
rect 35489 167023 35523 167051
rect 35551 167023 50697 167051
rect 50725 167023 50759 167051
rect 50787 167023 50821 167051
rect 50849 167023 50883 167051
rect 50911 167023 66057 167051
rect 66085 167023 66119 167051
rect 66147 167023 66181 167051
rect 66209 167023 66243 167051
rect 66271 167023 81417 167051
rect 81445 167023 81479 167051
rect 81507 167023 81541 167051
rect 81569 167023 81603 167051
rect 81631 167023 96777 167051
rect 96805 167023 96839 167051
rect 96867 167023 96901 167051
rect 96929 167023 96963 167051
rect 96991 167023 173577 167051
rect 173605 167023 173639 167051
rect 173667 167023 173701 167051
rect 173729 167023 173763 167051
rect 173791 167023 204297 167051
rect 204325 167023 204359 167051
rect 204387 167023 204421 167051
rect 204449 167023 204483 167051
rect 204511 167023 219657 167051
rect 219685 167023 219719 167051
rect 219747 167023 219781 167051
rect 219809 167023 219843 167051
rect 219871 167023 235017 167051
rect 235045 167023 235079 167051
rect 235107 167023 235141 167051
rect 235169 167023 235203 167051
rect 235231 167023 250377 167051
rect 250405 167023 250439 167051
rect 250467 167023 250501 167051
rect 250529 167023 250563 167051
rect 250591 167023 265737 167051
rect 265765 167023 265799 167051
rect 265827 167023 265861 167051
rect 265889 167023 265923 167051
rect 265951 167023 281097 167051
rect 281125 167023 281159 167051
rect 281187 167023 281221 167051
rect 281249 167023 281283 167051
rect 281311 167023 296457 167051
rect 296485 167023 296519 167051
rect 296547 167023 296581 167051
rect 296609 167023 296643 167051
rect 296671 167023 298728 167051
rect 298756 167023 298790 167051
rect 298818 167023 298852 167051
rect 298880 167023 298914 167051
rect 298942 167023 298990 167051
rect -958 166989 298990 167023
rect -958 166961 -910 166989
rect -882 166961 -848 166989
rect -820 166961 -786 166989
rect -758 166961 -724 166989
rect -696 166961 4617 166989
rect 4645 166961 4679 166989
rect 4707 166961 4741 166989
rect 4769 166961 4803 166989
rect 4831 166961 19977 166989
rect 20005 166961 20039 166989
rect 20067 166961 20101 166989
rect 20129 166961 20163 166989
rect 20191 166961 35337 166989
rect 35365 166961 35399 166989
rect 35427 166961 35461 166989
rect 35489 166961 35523 166989
rect 35551 166961 50697 166989
rect 50725 166961 50759 166989
rect 50787 166961 50821 166989
rect 50849 166961 50883 166989
rect 50911 166961 66057 166989
rect 66085 166961 66119 166989
rect 66147 166961 66181 166989
rect 66209 166961 66243 166989
rect 66271 166961 81417 166989
rect 81445 166961 81479 166989
rect 81507 166961 81541 166989
rect 81569 166961 81603 166989
rect 81631 166961 96777 166989
rect 96805 166961 96839 166989
rect 96867 166961 96901 166989
rect 96929 166961 96963 166989
rect 96991 166961 173577 166989
rect 173605 166961 173639 166989
rect 173667 166961 173701 166989
rect 173729 166961 173763 166989
rect 173791 166961 204297 166989
rect 204325 166961 204359 166989
rect 204387 166961 204421 166989
rect 204449 166961 204483 166989
rect 204511 166961 219657 166989
rect 219685 166961 219719 166989
rect 219747 166961 219781 166989
rect 219809 166961 219843 166989
rect 219871 166961 235017 166989
rect 235045 166961 235079 166989
rect 235107 166961 235141 166989
rect 235169 166961 235203 166989
rect 235231 166961 250377 166989
rect 250405 166961 250439 166989
rect 250467 166961 250501 166989
rect 250529 166961 250563 166989
rect 250591 166961 265737 166989
rect 265765 166961 265799 166989
rect 265827 166961 265861 166989
rect 265889 166961 265923 166989
rect 265951 166961 281097 166989
rect 281125 166961 281159 166989
rect 281187 166961 281221 166989
rect 281249 166961 281283 166989
rect 281311 166961 296457 166989
rect 296485 166961 296519 166989
rect 296547 166961 296581 166989
rect 296609 166961 296643 166989
rect 296671 166961 298728 166989
rect 298756 166961 298790 166989
rect 298818 166961 298852 166989
rect 298880 166961 298914 166989
rect 298942 166961 298990 166989
rect -958 166913 298990 166961
rect -958 164175 298990 164223
rect -958 164147 -430 164175
rect -402 164147 -368 164175
rect -340 164147 -306 164175
rect -278 164147 -244 164175
rect -216 164147 2757 164175
rect 2785 164147 2819 164175
rect 2847 164147 2881 164175
rect 2909 164147 2943 164175
rect 2971 164147 18117 164175
rect 18145 164147 18179 164175
rect 18207 164147 18241 164175
rect 18269 164147 18303 164175
rect 18331 164147 33477 164175
rect 33505 164147 33539 164175
rect 33567 164147 33601 164175
rect 33629 164147 33663 164175
rect 33691 164147 48837 164175
rect 48865 164147 48899 164175
rect 48927 164147 48961 164175
rect 48989 164147 49023 164175
rect 49051 164147 64197 164175
rect 64225 164147 64259 164175
rect 64287 164147 64321 164175
rect 64349 164147 64383 164175
rect 64411 164147 79557 164175
rect 79585 164147 79619 164175
rect 79647 164147 79681 164175
rect 79709 164147 79743 164175
rect 79771 164147 94917 164175
rect 94945 164147 94979 164175
rect 95007 164147 95041 164175
rect 95069 164147 95103 164175
rect 95131 164147 171717 164175
rect 171745 164147 171779 164175
rect 171807 164147 171841 164175
rect 171869 164147 171903 164175
rect 171931 164147 187077 164175
rect 187105 164147 187139 164175
rect 187167 164147 187201 164175
rect 187229 164147 187263 164175
rect 187291 164147 202437 164175
rect 202465 164147 202499 164175
rect 202527 164147 202561 164175
rect 202589 164147 202623 164175
rect 202651 164147 217797 164175
rect 217825 164147 217859 164175
rect 217887 164147 217921 164175
rect 217949 164147 217983 164175
rect 218011 164147 233157 164175
rect 233185 164147 233219 164175
rect 233247 164147 233281 164175
rect 233309 164147 233343 164175
rect 233371 164147 248517 164175
rect 248545 164147 248579 164175
rect 248607 164147 248641 164175
rect 248669 164147 248703 164175
rect 248731 164147 263877 164175
rect 263905 164147 263939 164175
rect 263967 164147 264001 164175
rect 264029 164147 264063 164175
rect 264091 164147 279237 164175
rect 279265 164147 279299 164175
rect 279327 164147 279361 164175
rect 279389 164147 279423 164175
rect 279451 164147 294597 164175
rect 294625 164147 294659 164175
rect 294687 164147 294721 164175
rect 294749 164147 294783 164175
rect 294811 164147 298248 164175
rect 298276 164147 298310 164175
rect 298338 164147 298372 164175
rect 298400 164147 298434 164175
rect 298462 164147 298990 164175
rect -958 164113 298990 164147
rect -958 164085 -430 164113
rect -402 164085 -368 164113
rect -340 164085 -306 164113
rect -278 164085 -244 164113
rect -216 164085 2757 164113
rect 2785 164085 2819 164113
rect 2847 164085 2881 164113
rect 2909 164085 2943 164113
rect 2971 164085 18117 164113
rect 18145 164085 18179 164113
rect 18207 164085 18241 164113
rect 18269 164085 18303 164113
rect 18331 164085 33477 164113
rect 33505 164085 33539 164113
rect 33567 164085 33601 164113
rect 33629 164085 33663 164113
rect 33691 164085 48837 164113
rect 48865 164085 48899 164113
rect 48927 164085 48961 164113
rect 48989 164085 49023 164113
rect 49051 164085 64197 164113
rect 64225 164085 64259 164113
rect 64287 164085 64321 164113
rect 64349 164085 64383 164113
rect 64411 164085 79557 164113
rect 79585 164085 79619 164113
rect 79647 164085 79681 164113
rect 79709 164085 79743 164113
rect 79771 164085 94917 164113
rect 94945 164085 94979 164113
rect 95007 164085 95041 164113
rect 95069 164085 95103 164113
rect 95131 164085 171717 164113
rect 171745 164085 171779 164113
rect 171807 164085 171841 164113
rect 171869 164085 171903 164113
rect 171931 164085 187077 164113
rect 187105 164085 187139 164113
rect 187167 164085 187201 164113
rect 187229 164085 187263 164113
rect 187291 164085 202437 164113
rect 202465 164085 202499 164113
rect 202527 164085 202561 164113
rect 202589 164085 202623 164113
rect 202651 164085 217797 164113
rect 217825 164085 217859 164113
rect 217887 164085 217921 164113
rect 217949 164085 217983 164113
rect 218011 164085 233157 164113
rect 233185 164085 233219 164113
rect 233247 164085 233281 164113
rect 233309 164085 233343 164113
rect 233371 164085 248517 164113
rect 248545 164085 248579 164113
rect 248607 164085 248641 164113
rect 248669 164085 248703 164113
rect 248731 164085 263877 164113
rect 263905 164085 263939 164113
rect 263967 164085 264001 164113
rect 264029 164085 264063 164113
rect 264091 164085 279237 164113
rect 279265 164085 279299 164113
rect 279327 164085 279361 164113
rect 279389 164085 279423 164113
rect 279451 164085 294597 164113
rect 294625 164085 294659 164113
rect 294687 164085 294721 164113
rect 294749 164085 294783 164113
rect 294811 164085 298248 164113
rect 298276 164085 298310 164113
rect 298338 164085 298372 164113
rect 298400 164085 298434 164113
rect 298462 164085 298990 164113
rect -958 164051 298990 164085
rect -958 164023 -430 164051
rect -402 164023 -368 164051
rect -340 164023 -306 164051
rect -278 164023 -244 164051
rect -216 164023 2757 164051
rect 2785 164023 2819 164051
rect 2847 164023 2881 164051
rect 2909 164023 2943 164051
rect 2971 164023 18117 164051
rect 18145 164023 18179 164051
rect 18207 164023 18241 164051
rect 18269 164023 18303 164051
rect 18331 164023 33477 164051
rect 33505 164023 33539 164051
rect 33567 164023 33601 164051
rect 33629 164023 33663 164051
rect 33691 164023 48837 164051
rect 48865 164023 48899 164051
rect 48927 164023 48961 164051
rect 48989 164023 49023 164051
rect 49051 164023 64197 164051
rect 64225 164023 64259 164051
rect 64287 164023 64321 164051
rect 64349 164023 64383 164051
rect 64411 164023 79557 164051
rect 79585 164023 79619 164051
rect 79647 164023 79681 164051
rect 79709 164023 79743 164051
rect 79771 164023 94917 164051
rect 94945 164023 94979 164051
rect 95007 164023 95041 164051
rect 95069 164023 95103 164051
rect 95131 164023 171717 164051
rect 171745 164023 171779 164051
rect 171807 164023 171841 164051
rect 171869 164023 171903 164051
rect 171931 164023 187077 164051
rect 187105 164023 187139 164051
rect 187167 164023 187201 164051
rect 187229 164023 187263 164051
rect 187291 164023 202437 164051
rect 202465 164023 202499 164051
rect 202527 164023 202561 164051
rect 202589 164023 202623 164051
rect 202651 164023 217797 164051
rect 217825 164023 217859 164051
rect 217887 164023 217921 164051
rect 217949 164023 217983 164051
rect 218011 164023 233157 164051
rect 233185 164023 233219 164051
rect 233247 164023 233281 164051
rect 233309 164023 233343 164051
rect 233371 164023 248517 164051
rect 248545 164023 248579 164051
rect 248607 164023 248641 164051
rect 248669 164023 248703 164051
rect 248731 164023 263877 164051
rect 263905 164023 263939 164051
rect 263967 164023 264001 164051
rect 264029 164023 264063 164051
rect 264091 164023 279237 164051
rect 279265 164023 279299 164051
rect 279327 164023 279361 164051
rect 279389 164023 279423 164051
rect 279451 164023 294597 164051
rect 294625 164023 294659 164051
rect 294687 164023 294721 164051
rect 294749 164023 294783 164051
rect 294811 164023 298248 164051
rect 298276 164023 298310 164051
rect 298338 164023 298372 164051
rect 298400 164023 298434 164051
rect 298462 164023 298990 164051
rect -958 163989 298990 164023
rect -958 163961 -430 163989
rect -402 163961 -368 163989
rect -340 163961 -306 163989
rect -278 163961 -244 163989
rect -216 163961 2757 163989
rect 2785 163961 2819 163989
rect 2847 163961 2881 163989
rect 2909 163961 2943 163989
rect 2971 163961 18117 163989
rect 18145 163961 18179 163989
rect 18207 163961 18241 163989
rect 18269 163961 18303 163989
rect 18331 163961 33477 163989
rect 33505 163961 33539 163989
rect 33567 163961 33601 163989
rect 33629 163961 33663 163989
rect 33691 163961 48837 163989
rect 48865 163961 48899 163989
rect 48927 163961 48961 163989
rect 48989 163961 49023 163989
rect 49051 163961 64197 163989
rect 64225 163961 64259 163989
rect 64287 163961 64321 163989
rect 64349 163961 64383 163989
rect 64411 163961 79557 163989
rect 79585 163961 79619 163989
rect 79647 163961 79681 163989
rect 79709 163961 79743 163989
rect 79771 163961 94917 163989
rect 94945 163961 94979 163989
rect 95007 163961 95041 163989
rect 95069 163961 95103 163989
rect 95131 163961 171717 163989
rect 171745 163961 171779 163989
rect 171807 163961 171841 163989
rect 171869 163961 171903 163989
rect 171931 163961 187077 163989
rect 187105 163961 187139 163989
rect 187167 163961 187201 163989
rect 187229 163961 187263 163989
rect 187291 163961 202437 163989
rect 202465 163961 202499 163989
rect 202527 163961 202561 163989
rect 202589 163961 202623 163989
rect 202651 163961 217797 163989
rect 217825 163961 217859 163989
rect 217887 163961 217921 163989
rect 217949 163961 217983 163989
rect 218011 163961 233157 163989
rect 233185 163961 233219 163989
rect 233247 163961 233281 163989
rect 233309 163961 233343 163989
rect 233371 163961 248517 163989
rect 248545 163961 248579 163989
rect 248607 163961 248641 163989
rect 248669 163961 248703 163989
rect 248731 163961 263877 163989
rect 263905 163961 263939 163989
rect 263967 163961 264001 163989
rect 264029 163961 264063 163989
rect 264091 163961 279237 163989
rect 279265 163961 279299 163989
rect 279327 163961 279361 163989
rect 279389 163961 279423 163989
rect 279451 163961 294597 163989
rect 294625 163961 294659 163989
rect 294687 163961 294721 163989
rect 294749 163961 294783 163989
rect 294811 163961 298248 163989
rect 298276 163961 298310 163989
rect 298338 163961 298372 163989
rect 298400 163961 298434 163989
rect 298462 163961 298990 163989
rect -958 163913 298990 163961
rect -958 158175 298990 158223
rect -958 158147 -910 158175
rect -882 158147 -848 158175
rect -820 158147 -786 158175
rect -758 158147 -724 158175
rect -696 158147 4617 158175
rect 4645 158147 4679 158175
rect 4707 158147 4741 158175
rect 4769 158147 4803 158175
rect 4831 158147 19977 158175
rect 20005 158147 20039 158175
rect 20067 158147 20101 158175
rect 20129 158147 20163 158175
rect 20191 158147 35337 158175
rect 35365 158147 35399 158175
rect 35427 158147 35461 158175
rect 35489 158147 35523 158175
rect 35551 158147 39939 158175
rect 39967 158147 40001 158175
rect 40029 158147 50697 158175
rect 50725 158147 50759 158175
rect 50787 158147 50821 158175
rect 50849 158147 50883 158175
rect 50911 158147 55299 158175
rect 55327 158147 55361 158175
rect 55389 158147 66057 158175
rect 66085 158147 66119 158175
rect 66147 158147 66181 158175
rect 66209 158147 66243 158175
rect 66271 158147 70659 158175
rect 70687 158147 70721 158175
rect 70749 158147 81417 158175
rect 81445 158147 81479 158175
rect 81507 158147 81541 158175
rect 81569 158147 81603 158175
rect 81631 158147 86019 158175
rect 86047 158147 86081 158175
rect 86109 158147 96777 158175
rect 96805 158147 96839 158175
rect 96867 158147 96901 158175
rect 96929 158147 96963 158175
rect 96991 158147 101379 158175
rect 101407 158147 101441 158175
rect 101469 158147 116739 158175
rect 116767 158147 116801 158175
rect 116829 158147 132099 158175
rect 132127 158147 132161 158175
rect 132189 158147 147459 158175
rect 147487 158147 147521 158175
rect 147549 158147 162819 158175
rect 162847 158147 162881 158175
rect 162909 158147 178179 158175
rect 178207 158147 178241 158175
rect 178269 158147 193539 158175
rect 193567 158147 193601 158175
rect 193629 158147 204297 158175
rect 204325 158147 204359 158175
rect 204387 158147 204421 158175
rect 204449 158147 204483 158175
rect 204511 158147 208899 158175
rect 208927 158147 208961 158175
rect 208989 158147 219657 158175
rect 219685 158147 219719 158175
rect 219747 158147 219781 158175
rect 219809 158147 219843 158175
rect 219871 158147 224259 158175
rect 224287 158147 224321 158175
rect 224349 158147 235017 158175
rect 235045 158147 235079 158175
rect 235107 158147 235141 158175
rect 235169 158147 235203 158175
rect 235231 158147 239619 158175
rect 239647 158147 239681 158175
rect 239709 158147 250377 158175
rect 250405 158147 250439 158175
rect 250467 158147 250501 158175
rect 250529 158147 250563 158175
rect 250591 158147 254979 158175
rect 255007 158147 255041 158175
rect 255069 158147 265737 158175
rect 265765 158147 265799 158175
rect 265827 158147 265861 158175
rect 265889 158147 265923 158175
rect 265951 158147 281097 158175
rect 281125 158147 281159 158175
rect 281187 158147 281221 158175
rect 281249 158147 281283 158175
rect 281311 158147 296457 158175
rect 296485 158147 296519 158175
rect 296547 158147 296581 158175
rect 296609 158147 296643 158175
rect 296671 158147 298728 158175
rect 298756 158147 298790 158175
rect 298818 158147 298852 158175
rect 298880 158147 298914 158175
rect 298942 158147 298990 158175
rect -958 158113 298990 158147
rect -958 158085 -910 158113
rect -882 158085 -848 158113
rect -820 158085 -786 158113
rect -758 158085 -724 158113
rect -696 158085 4617 158113
rect 4645 158085 4679 158113
rect 4707 158085 4741 158113
rect 4769 158085 4803 158113
rect 4831 158085 19977 158113
rect 20005 158085 20039 158113
rect 20067 158085 20101 158113
rect 20129 158085 20163 158113
rect 20191 158085 35337 158113
rect 35365 158085 35399 158113
rect 35427 158085 35461 158113
rect 35489 158085 35523 158113
rect 35551 158085 39939 158113
rect 39967 158085 40001 158113
rect 40029 158085 50697 158113
rect 50725 158085 50759 158113
rect 50787 158085 50821 158113
rect 50849 158085 50883 158113
rect 50911 158085 55299 158113
rect 55327 158085 55361 158113
rect 55389 158085 66057 158113
rect 66085 158085 66119 158113
rect 66147 158085 66181 158113
rect 66209 158085 66243 158113
rect 66271 158085 70659 158113
rect 70687 158085 70721 158113
rect 70749 158085 81417 158113
rect 81445 158085 81479 158113
rect 81507 158085 81541 158113
rect 81569 158085 81603 158113
rect 81631 158085 86019 158113
rect 86047 158085 86081 158113
rect 86109 158085 96777 158113
rect 96805 158085 96839 158113
rect 96867 158085 96901 158113
rect 96929 158085 96963 158113
rect 96991 158085 101379 158113
rect 101407 158085 101441 158113
rect 101469 158085 116739 158113
rect 116767 158085 116801 158113
rect 116829 158085 132099 158113
rect 132127 158085 132161 158113
rect 132189 158085 147459 158113
rect 147487 158085 147521 158113
rect 147549 158085 162819 158113
rect 162847 158085 162881 158113
rect 162909 158085 178179 158113
rect 178207 158085 178241 158113
rect 178269 158085 193539 158113
rect 193567 158085 193601 158113
rect 193629 158085 204297 158113
rect 204325 158085 204359 158113
rect 204387 158085 204421 158113
rect 204449 158085 204483 158113
rect 204511 158085 208899 158113
rect 208927 158085 208961 158113
rect 208989 158085 219657 158113
rect 219685 158085 219719 158113
rect 219747 158085 219781 158113
rect 219809 158085 219843 158113
rect 219871 158085 224259 158113
rect 224287 158085 224321 158113
rect 224349 158085 235017 158113
rect 235045 158085 235079 158113
rect 235107 158085 235141 158113
rect 235169 158085 235203 158113
rect 235231 158085 239619 158113
rect 239647 158085 239681 158113
rect 239709 158085 250377 158113
rect 250405 158085 250439 158113
rect 250467 158085 250501 158113
rect 250529 158085 250563 158113
rect 250591 158085 254979 158113
rect 255007 158085 255041 158113
rect 255069 158085 265737 158113
rect 265765 158085 265799 158113
rect 265827 158085 265861 158113
rect 265889 158085 265923 158113
rect 265951 158085 281097 158113
rect 281125 158085 281159 158113
rect 281187 158085 281221 158113
rect 281249 158085 281283 158113
rect 281311 158085 296457 158113
rect 296485 158085 296519 158113
rect 296547 158085 296581 158113
rect 296609 158085 296643 158113
rect 296671 158085 298728 158113
rect 298756 158085 298790 158113
rect 298818 158085 298852 158113
rect 298880 158085 298914 158113
rect 298942 158085 298990 158113
rect -958 158051 298990 158085
rect -958 158023 -910 158051
rect -882 158023 -848 158051
rect -820 158023 -786 158051
rect -758 158023 -724 158051
rect -696 158023 4617 158051
rect 4645 158023 4679 158051
rect 4707 158023 4741 158051
rect 4769 158023 4803 158051
rect 4831 158023 19977 158051
rect 20005 158023 20039 158051
rect 20067 158023 20101 158051
rect 20129 158023 20163 158051
rect 20191 158023 35337 158051
rect 35365 158023 35399 158051
rect 35427 158023 35461 158051
rect 35489 158023 35523 158051
rect 35551 158023 39939 158051
rect 39967 158023 40001 158051
rect 40029 158023 50697 158051
rect 50725 158023 50759 158051
rect 50787 158023 50821 158051
rect 50849 158023 50883 158051
rect 50911 158023 55299 158051
rect 55327 158023 55361 158051
rect 55389 158023 66057 158051
rect 66085 158023 66119 158051
rect 66147 158023 66181 158051
rect 66209 158023 66243 158051
rect 66271 158023 70659 158051
rect 70687 158023 70721 158051
rect 70749 158023 81417 158051
rect 81445 158023 81479 158051
rect 81507 158023 81541 158051
rect 81569 158023 81603 158051
rect 81631 158023 86019 158051
rect 86047 158023 86081 158051
rect 86109 158023 96777 158051
rect 96805 158023 96839 158051
rect 96867 158023 96901 158051
rect 96929 158023 96963 158051
rect 96991 158023 101379 158051
rect 101407 158023 101441 158051
rect 101469 158023 116739 158051
rect 116767 158023 116801 158051
rect 116829 158023 132099 158051
rect 132127 158023 132161 158051
rect 132189 158023 147459 158051
rect 147487 158023 147521 158051
rect 147549 158023 162819 158051
rect 162847 158023 162881 158051
rect 162909 158023 178179 158051
rect 178207 158023 178241 158051
rect 178269 158023 193539 158051
rect 193567 158023 193601 158051
rect 193629 158023 204297 158051
rect 204325 158023 204359 158051
rect 204387 158023 204421 158051
rect 204449 158023 204483 158051
rect 204511 158023 208899 158051
rect 208927 158023 208961 158051
rect 208989 158023 219657 158051
rect 219685 158023 219719 158051
rect 219747 158023 219781 158051
rect 219809 158023 219843 158051
rect 219871 158023 224259 158051
rect 224287 158023 224321 158051
rect 224349 158023 235017 158051
rect 235045 158023 235079 158051
rect 235107 158023 235141 158051
rect 235169 158023 235203 158051
rect 235231 158023 239619 158051
rect 239647 158023 239681 158051
rect 239709 158023 250377 158051
rect 250405 158023 250439 158051
rect 250467 158023 250501 158051
rect 250529 158023 250563 158051
rect 250591 158023 254979 158051
rect 255007 158023 255041 158051
rect 255069 158023 265737 158051
rect 265765 158023 265799 158051
rect 265827 158023 265861 158051
rect 265889 158023 265923 158051
rect 265951 158023 281097 158051
rect 281125 158023 281159 158051
rect 281187 158023 281221 158051
rect 281249 158023 281283 158051
rect 281311 158023 296457 158051
rect 296485 158023 296519 158051
rect 296547 158023 296581 158051
rect 296609 158023 296643 158051
rect 296671 158023 298728 158051
rect 298756 158023 298790 158051
rect 298818 158023 298852 158051
rect 298880 158023 298914 158051
rect 298942 158023 298990 158051
rect -958 157989 298990 158023
rect -958 157961 -910 157989
rect -882 157961 -848 157989
rect -820 157961 -786 157989
rect -758 157961 -724 157989
rect -696 157961 4617 157989
rect 4645 157961 4679 157989
rect 4707 157961 4741 157989
rect 4769 157961 4803 157989
rect 4831 157961 19977 157989
rect 20005 157961 20039 157989
rect 20067 157961 20101 157989
rect 20129 157961 20163 157989
rect 20191 157961 35337 157989
rect 35365 157961 35399 157989
rect 35427 157961 35461 157989
rect 35489 157961 35523 157989
rect 35551 157961 39939 157989
rect 39967 157961 40001 157989
rect 40029 157961 50697 157989
rect 50725 157961 50759 157989
rect 50787 157961 50821 157989
rect 50849 157961 50883 157989
rect 50911 157961 55299 157989
rect 55327 157961 55361 157989
rect 55389 157961 66057 157989
rect 66085 157961 66119 157989
rect 66147 157961 66181 157989
rect 66209 157961 66243 157989
rect 66271 157961 70659 157989
rect 70687 157961 70721 157989
rect 70749 157961 81417 157989
rect 81445 157961 81479 157989
rect 81507 157961 81541 157989
rect 81569 157961 81603 157989
rect 81631 157961 86019 157989
rect 86047 157961 86081 157989
rect 86109 157961 96777 157989
rect 96805 157961 96839 157989
rect 96867 157961 96901 157989
rect 96929 157961 96963 157989
rect 96991 157961 101379 157989
rect 101407 157961 101441 157989
rect 101469 157961 116739 157989
rect 116767 157961 116801 157989
rect 116829 157961 132099 157989
rect 132127 157961 132161 157989
rect 132189 157961 147459 157989
rect 147487 157961 147521 157989
rect 147549 157961 162819 157989
rect 162847 157961 162881 157989
rect 162909 157961 178179 157989
rect 178207 157961 178241 157989
rect 178269 157961 193539 157989
rect 193567 157961 193601 157989
rect 193629 157961 204297 157989
rect 204325 157961 204359 157989
rect 204387 157961 204421 157989
rect 204449 157961 204483 157989
rect 204511 157961 208899 157989
rect 208927 157961 208961 157989
rect 208989 157961 219657 157989
rect 219685 157961 219719 157989
rect 219747 157961 219781 157989
rect 219809 157961 219843 157989
rect 219871 157961 224259 157989
rect 224287 157961 224321 157989
rect 224349 157961 235017 157989
rect 235045 157961 235079 157989
rect 235107 157961 235141 157989
rect 235169 157961 235203 157989
rect 235231 157961 239619 157989
rect 239647 157961 239681 157989
rect 239709 157961 250377 157989
rect 250405 157961 250439 157989
rect 250467 157961 250501 157989
rect 250529 157961 250563 157989
rect 250591 157961 254979 157989
rect 255007 157961 255041 157989
rect 255069 157961 265737 157989
rect 265765 157961 265799 157989
rect 265827 157961 265861 157989
rect 265889 157961 265923 157989
rect 265951 157961 281097 157989
rect 281125 157961 281159 157989
rect 281187 157961 281221 157989
rect 281249 157961 281283 157989
rect 281311 157961 296457 157989
rect 296485 157961 296519 157989
rect 296547 157961 296581 157989
rect 296609 157961 296643 157989
rect 296671 157961 298728 157989
rect 298756 157961 298790 157989
rect 298818 157961 298852 157989
rect 298880 157961 298914 157989
rect 298942 157961 298990 157989
rect -958 157913 298990 157961
rect -958 155175 298990 155223
rect -958 155147 -430 155175
rect -402 155147 -368 155175
rect -340 155147 -306 155175
rect -278 155147 -244 155175
rect -216 155147 2757 155175
rect 2785 155147 2819 155175
rect 2847 155147 2881 155175
rect 2909 155147 2943 155175
rect 2971 155147 18117 155175
rect 18145 155147 18179 155175
rect 18207 155147 18241 155175
rect 18269 155147 18303 155175
rect 18331 155147 32259 155175
rect 32287 155147 32321 155175
rect 32349 155147 33477 155175
rect 33505 155147 33539 155175
rect 33567 155147 33601 155175
rect 33629 155147 33663 155175
rect 33691 155147 47619 155175
rect 47647 155147 47681 155175
rect 47709 155147 48837 155175
rect 48865 155147 48899 155175
rect 48927 155147 48961 155175
rect 48989 155147 49023 155175
rect 49051 155147 62979 155175
rect 63007 155147 63041 155175
rect 63069 155147 64197 155175
rect 64225 155147 64259 155175
rect 64287 155147 64321 155175
rect 64349 155147 64383 155175
rect 64411 155147 78339 155175
rect 78367 155147 78401 155175
rect 78429 155147 79557 155175
rect 79585 155147 79619 155175
rect 79647 155147 79681 155175
rect 79709 155147 79743 155175
rect 79771 155147 93699 155175
rect 93727 155147 93761 155175
rect 93789 155147 94917 155175
rect 94945 155147 94979 155175
rect 95007 155147 95041 155175
rect 95069 155147 95103 155175
rect 95131 155147 109059 155175
rect 109087 155147 109121 155175
rect 109149 155147 124419 155175
rect 124447 155147 124481 155175
rect 124509 155147 139779 155175
rect 139807 155147 139841 155175
rect 139869 155147 155139 155175
rect 155167 155147 155201 155175
rect 155229 155147 170499 155175
rect 170527 155147 170561 155175
rect 170589 155147 185859 155175
rect 185887 155147 185921 155175
rect 185949 155147 201219 155175
rect 201247 155147 201281 155175
rect 201309 155147 216579 155175
rect 216607 155147 216641 155175
rect 216669 155147 217797 155175
rect 217825 155147 217859 155175
rect 217887 155147 217921 155175
rect 217949 155147 217983 155175
rect 218011 155147 231939 155175
rect 231967 155147 232001 155175
rect 232029 155147 233157 155175
rect 233185 155147 233219 155175
rect 233247 155147 233281 155175
rect 233309 155147 233343 155175
rect 233371 155147 247299 155175
rect 247327 155147 247361 155175
rect 247389 155147 248517 155175
rect 248545 155147 248579 155175
rect 248607 155147 248641 155175
rect 248669 155147 248703 155175
rect 248731 155147 262659 155175
rect 262687 155147 262721 155175
rect 262749 155147 263877 155175
rect 263905 155147 263939 155175
rect 263967 155147 264001 155175
rect 264029 155147 264063 155175
rect 264091 155147 279237 155175
rect 279265 155147 279299 155175
rect 279327 155147 279361 155175
rect 279389 155147 279423 155175
rect 279451 155147 294597 155175
rect 294625 155147 294659 155175
rect 294687 155147 294721 155175
rect 294749 155147 294783 155175
rect 294811 155147 298248 155175
rect 298276 155147 298310 155175
rect 298338 155147 298372 155175
rect 298400 155147 298434 155175
rect 298462 155147 298990 155175
rect -958 155113 298990 155147
rect -958 155085 -430 155113
rect -402 155085 -368 155113
rect -340 155085 -306 155113
rect -278 155085 -244 155113
rect -216 155085 2757 155113
rect 2785 155085 2819 155113
rect 2847 155085 2881 155113
rect 2909 155085 2943 155113
rect 2971 155085 18117 155113
rect 18145 155085 18179 155113
rect 18207 155085 18241 155113
rect 18269 155085 18303 155113
rect 18331 155085 32259 155113
rect 32287 155085 32321 155113
rect 32349 155085 33477 155113
rect 33505 155085 33539 155113
rect 33567 155085 33601 155113
rect 33629 155085 33663 155113
rect 33691 155085 47619 155113
rect 47647 155085 47681 155113
rect 47709 155085 48837 155113
rect 48865 155085 48899 155113
rect 48927 155085 48961 155113
rect 48989 155085 49023 155113
rect 49051 155085 62979 155113
rect 63007 155085 63041 155113
rect 63069 155085 64197 155113
rect 64225 155085 64259 155113
rect 64287 155085 64321 155113
rect 64349 155085 64383 155113
rect 64411 155085 78339 155113
rect 78367 155085 78401 155113
rect 78429 155085 79557 155113
rect 79585 155085 79619 155113
rect 79647 155085 79681 155113
rect 79709 155085 79743 155113
rect 79771 155085 93699 155113
rect 93727 155085 93761 155113
rect 93789 155085 94917 155113
rect 94945 155085 94979 155113
rect 95007 155085 95041 155113
rect 95069 155085 95103 155113
rect 95131 155085 109059 155113
rect 109087 155085 109121 155113
rect 109149 155085 124419 155113
rect 124447 155085 124481 155113
rect 124509 155085 139779 155113
rect 139807 155085 139841 155113
rect 139869 155085 155139 155113
rect 155167 155085 155201 155113
rect 155229 155085 170499 155113
rect 170527 155085 170561 155113
rect 170589 155085 185859 155113
rect 185887 155085 185921 155113
rect 185949 155085 201219 155113
rect 201247 155085 201281 155113
rect 201309 155085 216579 155113
rect 216607 155085 216641 155113
rect 216669 155085 217797 155113
rect 217825 155085 217859 155113
rect 217887 155085 217921 155113
rect 217949 155085 217983 155113
rect 218011 155085 231939 155113
rect 231967 155085 232001 155113
rect 232029 155085 233157 155113
rect 233185 155085 233219 155113
rect 233247 155085 233281 155113
rect 233309 155085 233343 155113
rect 233371 155085 247299 155113
rect 247327 155085 247361 155113
rect 247389 155085 248517 155113
rect 248545 155085 248579 155113
rect 248607 155085 248641 155113
rect 248669 155085 248703 155113
rect 248731 155085 262659 155113
rect 262687 155085 262721 155113
rect 262749 155085 263877 155113
rect 263905 155085 263939 155113
rect 263967 155085 264001 155113
rect 264029 155085 264063 155113
rect 264091 155085 279237 155113
rect 279265 155085 279299 155113
rect 279327 155085 279361 155113
rect 279389 155085 279423 155113
rect 279451 155085 294597 155113
rect 294625 155085 294659 155113
rect 294687 155085 294721 155113
rect 294749 155085 294783 155113
rect 294811 155085 298248 155113
rect 298276 155085 298310 155113
rect 298338 155085 298372 155113
rect 298400 155085 298434 155113
rect 298462 155085 298990 155113
rect -958 155051 298990 155085
rect -958 155023 -430 155051
rect -402 155023 -368 155051
rect -340 155023 -306 155051
rect -278 155023 -244 155051
rect -216 155023 2757 155051
rect 2785 155023 2819 155051
rect 2847 155023 2881 155051
rect 2909 155023 2943 155051
rect 2971 155023 18117 155051
rect 18145 155023 18179 155051
rect 18207 155023 18241 155051
rect 18269 155023 18303 155051
rect 18331 155023 32259 155051
rect 32287 155023 32321 155051
rect 32349 155023 33477 155051
rect 33505 155023 33539 155051
rect 33567 155023 33601 155051
rect 33629 155023 33663 155051
rect 33691 155023 47619 155051
rect 47647 155023 47681 155051
rect 47709 155023 48837 155051
rect 48865 155023 48899 155051
rect 48927 155023 48961 155051
rect 48989 155023 49023 155051
rect 49051 155023 62979 155051
rect 63007 155023 63041 155051
rect 63069 155023 64197 155051
rect 64225 155023 64259 155051
rect 64287 155023 64321 155051
rect 64349 155023 64383 155051
rect 64411 155023 78339 155051
rect 78367 155023 78401 155051
rect 78429 155023 79557 155051
rect 79585 155023 79619 155051
rect 79647 155023 79681 155051
rect 79709 155023 79743 155051
rect 79771 155023 93699 155051
rect 93727 155023 93761 155051
rect 93789 155023 94917 155051
rect 94945 155023 94979 155051
rect 95007 155023 95041 155051
rect 95069 155023 95103 155051
rect 95131 155023 109059 155051
rect 109087 155023 109121 155051
rect 109149 155023 124419 155051
rect 124447 155023 124481 155051
rect 124509 155023 139779 155051
rect 139807 155023 139841 155051
rect 139869 155023 155139 155051
rect 155167 155023 155201 155051
rect 155229 155023 170499 155051
rect 170527 155023 170561 155051
rect 170589 155023 185859 155051
rect 185887 155023 185921 155051
rect 185949 155023 201219 155051
rect 201247 155023 201281 155051
rect 201309 155023 216579 155051
rect 216607 155023 216641 155051
rect 216669 155023 217797 155051
rect 217825 155023 217859 155051
rect 217887 155023 217921 155051
rect 217949 155023 217983 155051
rect 218011 155023 231939 155051
rect 231967 155023 232001 155051
rect 232029 155023 233157 155051
rect 233185 155023 233219 155051
rect 233247 155023 233281 155051
rect 233309 155023 233343 155051
rect 233371 155023 247299 155051
rect 247327 155023 247361 155051
rect 247389 155023 248517 155051
rect 248545 155023 248579 155051
rect 248607 155023 248641 155051
rect 248669 155023 248703 155051
rect 248731 155023 262659 155051
rect 262687 155023 262721 155051
rect 262749 155023 263877 155051
rect 263905 155023 263939 155051
rect 263967 155023 264001 155051
rect 264029 155023 264063 155051
rect 264091 155023 279237 155051
rect 279265 155023 279299 155051
rect 279327 155023 279361 155051
rect 279389 155023 279423 155051
rect 279451 155023 294597 155051
rect 294625 155023 294659 155051
rect 294687 155023 294721 155051
rect 294749 155023 294783 155051
rect 294811 155023 298248 155051
rect 298276 155023 298310 155051
rect 298338 155023 298372 155051
rect 298400 155023 298434 155051
rect 298462 155023 298990 155051
rect -958 154989 298990 155023
rect -958 154961 -430 154989
rect -402 154961 -368 154989
rect -340 154961 -306 154989
rect -278 154961 -244 154989
rect -216 154961 2757 154989
rect 2785 154961 2819 154989
rect 2847 154961 2881 154989
rect 2909 154961 2943 154989
rect 2971 154961 18117 154989
rect 18145 154961 18179 154989
rect 18207 154961 18241 154989
rect 18269 154961 18303 154989
rect 18331 154961 32259 154989
rect 32287 154961 32321 154989
rect 32349 154961 33477 154989
rect 33505 154961 33539 154989
rect 33567 154961 33601 154989
rect 33629 154961 33663 154989
rect 33691 154961 47619 154989
rect 47647 154961 47681 154989
rect 47709 154961 48837 154989
rect 48865 154961 48899 154989
rect 48927 154961 48961 154989
rect 48989 154961 49023 154989
rect 49051 154961 62979 154989
rect 63007 154961 63041 154989
rect 63069 154961 64197 154989
rect 64225 154961 64259 154989
rect 64287 154961 64321 154989
rect 64349 154961 64383 154989
rect 64411 154961 78339 154989
rect 78367 154961 78401 154989
rect 78429 154961 79557 154989
rect 79585 154961 79619 154989
rect 79647 154961 79681 154989
rect 79709 154961 79743 154989
rect 79771 154961 93699 154989
rect 93727 154961 93761 154989
rect 93789 154961 94917 154989
rect 94945 154961 94979 154989
rect 95007 154961 95041 154989
rect 95069 154961 95103 154989
rect 95131 154961 109059 154989
rect 109087 154961 109121 154989
rect 109149 154961 124419 154989
rect 124447 154961 124481 154989
rect 124509 154961 139779 154989
rect 139807 154961 139841 154989
rect 139869 154961 155139 154989
rect 155167 154961 155201 154989
rect 155229 154961 170499 154989
rect 170527 154961 170561 154989
rect 170589 154961 185859 154989
rect 185887 154961 185921 154989
rect 185949 154961 201219 154989
rect 201247 154961 201281 154989
rect 201309 154961 216579 154989
rect 216607 154961 216641 154989
rect 216669 154961 217797 154989
rect 217825 154961 217859 154989
rect 217887 154961 217921 154989
rect 217949 154961 217983 154989
rect 218011 154961 231939 154989
rect 231967 154961 232001 154989
rect 232029 154961 233157 154989
rect 233185 154961 233219 154989
rect 233247 154961 233281 154989
rect 233309 154961 233343 154989
rect 233371 154961 247299 154989
rect 247327 154961 247361 154989
rect 247389 154961 248517 154989
rect 248545 154961 248579 154989
rect 248607 154961 248641 154989
rect 248669 154961 248703 154989
rect 248731 154961 262659 154989
rect 262687 154961 262721 154989
rect 262749 154961 263877 154989
rect 263905 154961 263939 154989
rect 263967 154961 264001 154989
rect 264029 154961 264063 154989
rect 264091 154961 279237 154989
rect 279265 154961 279299 154989
rect 279327 154961 279361 154989
rect 279389 154961 279423 154989
rect 279451 154961 294597 154989
rect 294625 154961 294659 154989
rect 294687 154961 294721 154989
rect 294749 154961 294783 154989
rect 294811 154961 298248 154989
rect 298276 154961 298310 154989
rect 298338 154961 298372 154989
rect 298400 154961 298434 154989
rect 298462 154961 298990 154989
rect -958 154913 298990 154961
rect -958 149175 298990 149223
rect -958 149147 -910 149175
rect -882 149147 -848 149175
rect -820 149147 -786 149175
rect -758 149147 -724 149175
rect -696 149147 4617 149175
rect 4645 149147 4679 149175
rect 4707 149147 4741 149175
rect 4769 149147 4803 149175
rect 4831 149147 19977 149175
rect 20005 149147 20039 149175
rect 20067 149147 20101 149175
rect 20129 149147 20163 149175
rect 20191 149147 35337 149175
rect 35365 149147 35399 149175
rect 35427 149147 35461 149175
rect 35489 149147 35523 149175
rect 35551 149147 39939 149175
rect 39967 149147 40001 149175
rect 40029 149147 50697 149175
rect 50725 149147 50759 149175
rect 50787 149147 50821 149175
rect 50849 149147 50883 149175
rect 50911 149147 55299 149175
rect 55327 149147 55361 149175
rect 55389 149147 66057 149175
rect 66085 149147 66119 149175
rect 66147 149147 66181 149175
rect 66209 149147 66243 149175
rect 66271 149147 70659 149175
rect 70687 149147 70721 149175
rect 70749 149147 81417 149175
rect 81445 149147 81479 149175
rect 81507 149147 81541 149175
rect 81569 149147 81603 149175
rect 81631 149147 86019 149175
rect 86047 149147 86081 149175
rect 86109 149147 96777 149175
rect 96805 149147 96839 149175
rect 96867 149147 96901 149175
rect 96929 149147 96963 149175
rect 96991 149147 101379 149175
rect 101407 149147 101441 149175
rect 101469 149147 116739 149175
rect 116767 149147 116801 149175
rect 116829 149147 132099 149175
rect 132127 149147 132161 149175
rect 132189 149147 147459 149175
rect 147487 149147 147521 149175
rect 147549 149147 162819 149175
rect 162847 149147 162881 149175
rect 162909 149147 178179 149175
rect 178207 149147 178241 149175
rect 178269 149147 193539 149175
rect 193567 149147 193601 149175
rect 193629 149147 204297 149175
rect 204325 149147 204359 149175
rect 204387 149147 204421 149175
rect 204449 149147 204483 149175
rect 204511 149147 208899 149175
rect 208927 149147 208961 149175
rect 208989 149147 219657 149175
rect 219685 149147 219719 149175
rect 219747 149147 219781 149175
rect 219809 149147 219843 149175
rect 219871 149147 224259 149175
rect 224287 149147 224321 149175
rect 224349 149147 235017 149175
rect 235045 149147 235079 149175
rect 235107 149147 235141 149175
rect 235169 149147 235203 149175
rect 235231 149147 239619 149175
rect 239647 149147 239681 149175
rect 239709 149147 250377 149175
rect 250405 149147 250439 149175
rect 250467 149147 250501 149175
rect 250529 149147 250563 149175
rect 250591 149147 254979 149175
rect 255007 149147 255041 149175
rect 255069 149147 265737 149175
rect 265765 149147 265799 149175
rect 265827 149147 265861 149175
rect 265889 149147 265923 149175
rect 265951 149147 281097 149175
rect 281125 149147 281159 149175
rect 281187 149147 281221 149175
rect 281249 149147 281283 149175
rect 281311 149147 296457 149175
rect 296485 149147 296519 149175
rect 296547 149147 296581 149175
rect 296609 149147 296643 149175
rect 296671 149147 298728 149175
rect 298756 149147 298790 149175
rect 298818 149147 298852 149175
rect 298880 149147 298914 149175
rect 298942 149147 298990 149175
rect -958 149113 298990 149147
rect -958 149085 -910 149113
rect -882 149085 -848 149113
rect -820 149085 -786 149113
rect -758 149085 -724 149113
rect -696 149085 4617 149113
rect 4645 149085 4679 149113
rect 4707 149085 4741 149113
rect 4769 149085 4803 149113
rect 4831 149085 19977 149113
rect 20005 149085 20039 149113
rect 20067 149085 20101 149113
rect 20129 149085 20163 149113
rect 20191 149085 35337 149113
rect 35365 149085 35399 149113
rect 35427 149085 35461 149113
rect 35489 149085 35523 149113
rect 35551 149085 39939 149113
rect 39967 149085 40001 149113
rect 40029 149085 50697 149113
rect 50725 149085 50759 149113
rect 50787 149085 50821 149113
rect 50849 149085 50883 149113
rect 50911 149085 55299 149113
rect 55327 149085 55361 149113
rect 55389 149085 66057 149113
rect 66085 149085 66119 149113
rect 66147 149085 66181 149113
rect 66209 149085 66243 149113
rect 66271 149085 70659 149113
rect 70687 149085 70721 149113
rect 70749 149085 81417 149113
rect 81445 149085 81479 149113
rect 81507 149085 81541 149113
rect 81569 149085 81603 149113
rect 81631 149085 86019 149113
rect 86047 149085 86081 149113
rect 86109 149085 96777 149113
rect 96805 149085 96839 149113
rect 96867 149085 96901 149113
rect 96929 149085 96963 149113
rect 96991 149085 101379 149113
rect 101407 149085 101441 149113
rect 101469 149085 116739 149113
rect 116767 149085 116801 149113
rect 116829 149085 132099 149113
rect 132127 149085 132161 149113
rect 132189 149085 147459 149113
rect 147487 149085 147521 149113
rect 147549 149085 162819 149113
rect 162847 149085 162881 149113
rect 162909 149085 178179 149113
rect 178207 149085 178241 149113
rect 178269 149085 193539 149113
rect 193567 149085 193601 149113
rect 193629 149085 204297 149113
rect 204325 149085 204359 149113
rect 204387 149085 204421 149113
rect 204449 149085 204483 149113
rect 204511 149085 208899 149113
rect 208927 149085 208961 149113
rect 208989 149085 219657 149113
rect 219685 149085 219719 149113
rect 219747 149085 219781 149113
rect 219809 149085 219843 149113
rect 219871 149085 224259 149113
rect 224287 149085 224321 149113
rect 224349 149085 235017 149113
rect 235045 149085 235079 149113
rect 235107 149085 235141 149113
rect 235169 149085 235203 149113
rect 235231 149085 239619 149113
rect 239647 149085 239681 149113
rect 239709 149085 250377 149113
rect 250405 149085 250439 149113
rect 250467 149085 250501 149113
rect 250529 149085 250563 149113
rect 250591 149085 254979 149113
rect 255007 149085 255041 149113
rect 255069 149085 265737 149113
rect 265765 149085 265799 149113
rect 265827 149085 265861 149113
rect 265889 149085 265923 149113
rect 265951 149085 281097 149113
rect 281125 149085 281159 149113
rect 281187 149085 281221 149113
rect 281249 149085 281283 149113
rect 281311 149085 296457 149113
rect 296485 149085 296519 149113
rect 296547 149085 296581 149113
rect 296609 149085 296643 149113
rect 296671 149085 298728 149113
rect 298756 149085 298790 149113
rect 298818 149085 298852 149113
rect 298880 149085 298914 149113
rect 298942 149085 298990 149113
rect -958 149051 298990 149085
rect -958 149023 -910 149051
rect -882 149023 -848 149051
rect -820 149023 -786 149051
rect -758 149023 -724 149051
rect -696 149023 4617 149051
rect 4645 149023 4679 149051
rect 4707 149023 4741 149051
rect 4769 149023 4803 149051
rect 4831 149023 19977 149051
rect 20005 149023 20039 149051
rect 20067 149023 20101 149051
rect 20129 149023 20163 149051
rect 20191 149023 35337 149051
rect 35365 149023 35399 149051
rect 35427 149023 35461 149051
rect 35489 149023 35523 149051
rect 35551 149023 39939 149051
rect 39967 149023 40001 149051
rect 40029 149023 50697 149051
rect 50725 149023 50759 149051
rect 50787 149023 50821 149051
rect 50849 149023 50883 149051
rect 50911 149023 55299 149051
rect 55327 149023 55361 149051
rect 55389 149023 66057 149051
rect 66085 149023 66119 149051
rect 66147 149023 66181 149051
rect 66209 149023 66243 149051
rect 66271 149023 70659 149051
rect 70687 149023 70721 149051
rect 70749 149023 81417 149051
rect 81445 149023 81479 149051
rect 81507 149023 81541 149051
rect 81569 149023 81603 149051
rect 81631 149023 86019 149051
rect 86047 149023 86081 149051
rect 86109 149023 96777 149051
rect 96805 149023 96839 149051
rect 96867 149023 96901 149051
rect 96929 149023 96963 149051
rect 96991 149023 101379 149051
rect 101407 149023 101441 149051
rect 101469 149023 116739 149051
rect 116767 149023 116801 149051
rect 116829 149023 132099 149051
rect 132127 149023 132161 149051
rect 132189 149023 147459 149051
rect 147487 149023 147521 149051
rect 147549 149023 162819 149051
rect 162847 149023 162881 149051
rect 162909 149023 178179 149051
rect 178207 149023 178241 149051
rect 178269 149023 193539 149051
rect 193567 149023 193601 149051
rect 193629 149023 204297 149051
rect 204325 149023 204359 149051
rect 204387 149023 204421 149051
rect 204449 149023 204483 149051
rect 204511 149023 208899 149051
rect 208927 149023 208961 149051
rect 208989 149023 219657 149051
rect 219685 149023 219719 149051
rect 219747 149023 219781 149051
rect 219809 149023 219843 149051
rect 219871 149023 224259 149051
rect 224287 149023 224321 149051
rect 224349 149023 235017 149051
rect 235045 149023 235079 149051
rect 235107 149023 235141 149051
rect 235169 149023 235203 149051
rect 235231 149023 239619 149051
rect 239647 149023 239681 149051
rect 239709 149023 250377 149051
rect 250405 149023 250439 149051
rect 250467 149023 250501 149051
rect 250529 149023 250563 149051
rect 250591 149023 254979 149051
rect 255007 149023 255041 149051
rect 255069 149023 265737 149051
rect 265765 149023 265799 149051
rect 265827 149023 265861 149051
rect 265889 149023 265923 149051
rect 265951 149023 281097 149051
rect 281125 149023 281159 149051
rect 281187 149023 281221 149051
rect 281249 149023 281283 149051
rect 281311 149023 296457 149051
rect 296485 149023 296519 149051
rect 296547 149023 296581 149051
rect 296609 149023 296643 149051
rect 296671 149023 298728 149051
rect 298756 149023 298790 149051
rect 298818 149023 298852 149051
rect 298880 149023 298914 149051
rect 298942 149023 298990 149051
rect -958 148989 298990 149023
rect -958 148961 -910 148989
rect -882 148961 -848 148989
rect -820 148961 -786 148989
rect -758 148961 -724 148989
rect -696 148961 4617 148989
rect 4645 148961 4679 148989
rect 4707 148961 4741 148989
rect 4769 148961 4803 148989
rect 4831 148961 19977 148989
rect 20005 148961 20039 148989
rect 20067 148961 20101 148989
rect 20129 148961 20163 148989
rect 20191 148961 35337 148989
rect 35365 148961 35399 148989
rect 35427 148961 35461 148989
rect 35489 148961 35523 148989
rect 35551 148961 39939 148989
rect 39967 148961 40001 148989
rect 40029 148961 50697 148989
rect 50725 148961 50759 148989
rect 50787 148961 50821 148989
rect 50849 148961 50883 148989
rect 50911 148961 55299 148989
rect 55327 148961 55361 148989
rect 55389 148961 66057 148989
rect 66085 148961 66119 148989
rect 66147 148961 66181 148989
rect 66209 148961 66243 148989
rect 66271 148961 70659 148989
rect 70687 148961 70721 148989
rect 70749 148961 81417 148989
rect 81445 148961 81479 148989
rect 81507 148961 81541 148989
rect 81569 148961 81603 148989
rect 81631 148961 86019 148989
rect 86047 148961 86081 148989
rect 86109 148961 96777 148989
rect 96805 148961 96839 148989
rect 96867 148961 96901 148989
rect 96929 148961 96963 148989
rect 96991 148961 101379 148989
rect 101407 148961 101441 148989
rect 101469 148961 116739 148989
rect 116767 148961 116801 148989
rect 116829 148961 132099 148989
rect 132127 148961 132161 148989
rect 132189 148961 147459 148989
rect 147487 148961 147521 148989
rect 147549 148961 162819 148989
rect 162847 148961 162881 148989
rect 162909 148961 178179 148989
rect 178207 148961 178241 148989
rect 178269 148961 193539 148989
rect 193567 148961 193601 148989
rect 193629 148961 204297 148989
rect 204325 148961 204359 148989
rect 204387 148961 204421 148989
rect 204449 148961 204483 148989
rect 204511 148961 208899 148989
rect 208927 148961 208961 148989
rect 208989 148961 219657 148989
rect 219685 148961 219719 148989
rect 219747 148961 219781 148989
rect 219809 148961 219843 148989
rect 219871 148961 224259 148989
rect 224287 148961 224321 148989
rect 224349 148961 235017 148989
rect 235045 148961 235079 148989
rect 235107 148961 235141 148989
rect 235169 148961 235203 148989
rect 235231 148961 239619 148989
rect 239647 148961 239681 148989
rect 239709 148961 250377 148989
rect 250405 148961 250439 148989
rect 250467 148961 250501 148989
rect 250529 148961 250563 148989
rect 250591 148961 254979 148989
rect 255007 148961 255041 148989
rect 255069 148961 265737 148989
rect 265765 148961 265799 148989
rect 265827 148961 265861 148989
rect 265889 148961 265923 148989
rect 265951 148961 281097 148989
rect 281125 148961 281159 148989
rect 281187 148961 281221 148989
rect 281249 148961 281283 148989
rect 281311 148961 296457 148989
rect 296485 148961 296519 148989
rect 296547 148961 296581 148989
rect 296609 148961 296643 148989
rect 296671 148961 298728 148989
rect 298756 148961 298790 148989
rect 298818 148961 298852 148989
rect 298880 148961 298914 148989
rect 298942 148961 298990 148989
rect -958 148913 298990 148961
rect -958 146175 298990 146223
rect -958 146147 -430 146175
rect -402 146147 -368 146175
rect -340 146147 -306 146175
rect -278 146147 -244 146175
rect -216 146147 2757 146175
rect 2785 146147 2819 146175
rect 2847 146147 2881 146175
rect 2909 146147 2943 146175
rect 2971 146147 18117 146175
rect 18145 146147 18179 146175
rect 18207 146147 18241 146175
rect 18269 146147 18303 146175
rect 18331 146147 32259 146175
rect 32287 146147 32321 146175
rect 32349 146147 33477 146175
rect 33505 146147 33539 146175
rect 33567 146147 33601 146175
rect 33629 146147 33663 146175
rect 33691 146147 47619 146175
rect 47647 146147 47681 146175
rect 47709 146147 48837 146175
rect 48865 146147 48899 146175
rect 48927 146147 48961 146175
rect 48989 146147 49023 146175
rect 49051 146147 62979 146175
rect 63007 146147 63041 146175
rect 63069 146147 64197 146175
rect 64225 146147 64259 146175
rect 64287 146147 64321 146175
rect 64349 146147 64383 146175
rect 64411 146147 78339 146175
rect 78367 146147 78401 146175
rect 78429 146147 79557 146175
rect 79585 146147 79619 146175
rect 79647 146147 79681 146175
rect 79709 146147 79743 146175
rect 79771 146147 93699 146175
rect 93727 146147 93761 146175
rect 93789 146147 94917 146175
rect 94945 146147 94979 146175
rect 95007 146147 95041 146175
rect 95069 146147 95103 146175
rect 95131 146147 109059 146175
rect 109087 146147 109121 146175
rect 109149 146147 124419 146175
rect 124447 146147 124481 146175
rect 124509 146147 139779 146175
rect 139807 146147 139841 146175
rect 139869 146147 155139 146175
rect 155167 146147 155201 146175
rect 155229 146147 170499 146175
rect 170527 146147 170561 146175
rect 170589 146147 185859 146175
rect 185887 146147 185921 146175
rect 185949 146147 201219 146175
rect 201247 146147 201281 146175
rect 201309 146147 216579 146175
rect 216607 146147 216641 146175
rect 216669 146147 217797 146175
rect 217825 146147 217859 146175
rect 217887 146147 217921 146175
rect 217949 146147 217983 146175
rect 218011 146147 231939 146175
rect 231967 146147 232001 146175
rect 232029 146147 233157 146175
rect 233185 146147 233219 146175
rect 233247 146147 233281 146175
rect 233309 146147 233343 146175
rect 233371 146147 247299 146175
rect 247327 146147 247361 146175
rect 247389 146147 248517 146175
rect 248545 146147 248579 146175
rect 248607 146147 248641 146175
rect 248669 146147 248703 146175
rect 248731 146147 262659 146175
rect 262687 146147 262721 146175
rect 262749 146147 263877 146175
rect 263905 146147 263939 146175
rect 263967 146147 264001 146175
rect 264029 146147 264063 146175
rect 264091 146147 279237 146175
rect 279265 146147 279299 146175
rect 279327 146147 279361 146175
rect 279389 146147 279423 146175
rect 279451 146147 294597 146175
rect 294625 146147 294659 146175
rect 294687 146147 294721 146175
rect 294749 146147 294783 146175
rect 294811 146147 298248 146175
rect 298276 146147 298310 146175
rect 298338 146147 298372 146175
rect 298400 146147 298434 146175
rect 298462 146147 298990 146175
rect -958 146113 298990 146147
rect -958 146085 -430 146113
rect -402 146085 -368 146113
rect -340 146085 -306 146113
rect -278 146085 -244 146113
rect -216 146085 2757 146113
rect 2785 146085 2819 146113
rect 2847 146085 2881 146113
rect 2909 146085 2943 146113
rect 2971 146085 18117 146113
rect 18145 146085 18179 146113
rect 18207 146085 18241 146113
rect 18269 146085 18303 146113
rect 18331 146085 32259 146113
rect 32287 146085 32321 146113
rect 32349 146085 33477 146113
rect 33505 146085 33539 146113
rect 33567 146085 33601 146113
rect 33629 146085 33663 146113
rect 33691 146085 47619 146113
rect 47647 146085 47681 146113
rect 47709 146085 48837 146113
rect 48865 146085 48899 146113
rect 48927 146085 48961 146113
rect 48989 146085 49023 146113
rect 49051 146085 62979 146113
rect 63007 146085 63041 146113
rect 63069 146085 64197 146113
rect 64225 146085 64259 146113
rect 64287 146085 64321 146113
rect 64349 146085 64383 146113
rect 64411 146085 78339 146113
rect 78367 146085 78401 146113
rect 78429 146085 79557 146113
rect 79585 146085 79619 146113
rect 79647 146085 79681 146113
rect 79709 146085 79743 146113
rect 79771 146085 93699 146113
rect 93727 146085 93761 146113
rect 93789 146085 94917 146113
rect 94945 146085 94979 146113
rect 95007 146085 95041 146113
rect 95069 146085 95103 146113
rect 95131 146085 109059 146113
rect 109087 146085 109121 146113
rect 109149 146085 124419 146113
rect 124447 146085 124481 146113
rect 124509 146085 139779 146113
rect 139807 146085 139841 146113
rect 139869 146085 155139 146113
rect 155167 146085 155201 146113
rect 155229 146085 170499 146113
rect 170527 146085 170561 146113
rect 170589 146085 185859 146113
rect 185887 146085 185921 146113
rect 185949 146085 201219 146113
rect 201247 146085 201281 146113
rect 201309 146085 216579 146113
rect 216607 146085 216641 146113
rect 216669 146085 217797 146113
rect 217825 146085 217859 146113
rect 217887 146085 217921 146113
rect 217949 146085 217983 146113
rect 218011 146085 231939 146113
rect 231967 146085 232001 146113
rect 232029 146085 233157 146113
rect 233185 146085 233219 146113
rect 233247 146085 233281 146113
rect 233309 146085 233343 146113
rect 233371 146085 247299 146113
rect 247327 146085 247361 146113
rect 247389 146085 248517 146113
rect 248545 146085 248579 146113
rect 248607 146085 248641 146113
rect 248669 146085 248703 146113
rect 248731 146085 262659 146113
rect 262687 146085 262721 146113
rect 262749 146085 263877 146113
rect 263905 146085 263939 146113
rect 263967 146085 264001 146113
rect 264029 146085 264063 146113
rect 264091 146085 279237 146113
rect 279265 146085 279299 146113
rect 279327 146085 279361 146113
rect 279389 146085 279423 146113
rect 279451 146085 294597 146113
rect 294625 146085 294659 146113
rect 294687 146085 294721 146113
rect 294749 146085 294783 146113
rect 294811 146085 298248 146113
rect 298276 146085 298310 146113
rect 298338 146085 298372 146113
rect 298400 146085 298434 146113
rect 298462 146085 298990 146113
rect -958 146051 298990 146085
rect -958 146023 -430 146051
rect -402 146023 -368 146051
rect -340 146023 -306 146051
rect -278 146023 -244 146051
rect -216 146023 2757 146051
rect 2785 146023 2819 146051
rect 2847 146023 2881 146051
rect 2909 146023 2943 146051
rect 2971 146023 18117 146051
rect 18145 146023 18179 146051
rect 18207 146023 18241 146051
rect 18269 146023 18303 146051
rect 18331 146023 32259 146051
rect 32287 146023 32321 146051
rect 32349 146023 33477 146051
rect 33505 146023 33539 146051
rect 33567 146023 33601 146051
rect 33629 146023 33663 146051
rect 33691 146023 47619 146051
rect 47647 146023 47681 146051
rect 47709 146023 48837 146051
rect 48865 146023 48899 146051
rect 48927 146023 48961 146051
rect 48989 146023 49023 146051
rect 49051 146023 62979 146051
rect 63007 146023 63041 146051
rect 63069 146023 64197 146051
rect 64225 146023 64259 146051
rect 64287 146023 64321 146051
rect 64349 146023 64383 146051
rect 64411 146023 78339 146051
rect 78367 146023 78401 146051
rect 78429 146023 79557 146051
rect 79585 146023 79619 146051
rect 79647 146023 79681 146051
rect 79709 146023 79743 146051
rect 79771 146023 93699 146051
rect 93727 146023 93761 146051
rect 93789 146023 94917 146051
rect 94945 146023 94979 146051
rect 95007 146023 95041 146051
rect 95069 146023 95103 146051
rect 95131 146023 109059 146051
rect 109087 146023 109121 146051
rect 109149 146023 124419 146051
rect 124447 146023 124481 146051
rect 124509 146023 139779 146051
rect 139807 146023 139841 146051
rect 139869 146023 155139 146051
rect 155167 146023 155201 146051
rect 155229 146023 170499 146051
rect 170527 146023 170561 146051
rect 170589 146023 185859 146051
rect 185887 146023 185921 146051
rect 185949 146023 201219 146051
rect 201247 146023 201281 146051
rect 201309 146023 216579 146051
rect 216607 146023 216641 146051
rect 216669 146023 217797 146051
rect 217825 146023 217859 146051
rect 217887 146023 217921 146051
rect 217949 146023 217983 146051
rect 218011 146023 231939 146051
rect 231967 146023 232001 146051
rect 232029 146023 233157 146051
rect 233185 146023 233219 146051
rect 233247 146023 233281 146051
rect 233309 146023 233343 146051
rect 233371 146023 247299 146051
rect 247327 146023 247361 146051
rect 247389 146023 248517 146051
rect 248545 146023 248579 146051
rect 248607 146023 248641 146051
rect 248669 146023 248703 146051
rect 248731 146023 262659 146051
rect 262687 146023 262721 146051
rect 262749 146023 263877 146051
rect 263905 146023 263939 146051
rect 263967 146023 264001 146051
rect 264029 146023 264063 146051
rect 264091 146023 279237 146051
rect 279265 146023 279299 146051
rect 279327 146023 279361 146051
rect 279389 146023 279423 146051
rect 279451 146023 294597 146051
rect 294625 146023 294659 146051
rect 294687 146023 294721 146051
rect 294749 146023 294783 146051
rect 294811 146023 298248 146051
rect 298276 146023 298310 146051
rect 298338 146023 298372 146051
rect 298400 146023 298434 146051
rect 298462 146023 298990 146051
rect -958 145989 298990 146023
rect -958 145961 -430 145989
rect -402 145961 -368 145989
rect -340 145961 -306 145989
rect -278 145961 -244 145989
rect -216 145961 2757 145989
rect 2785 145961 2819 145989
rect 2847 145961 2881 145989
rect 2909 145961 2943 145989
rect 2971 145961 18117 145989
rect 18145 145961 18179 145989
rect 18207 145961 18241 145989
rect 18269 145961 18303 145989
rect 18331 145961 32259 145989
rect 32287 145961 32321 145989
rect 32349 145961 33477 145989
rect 33505 145961 33539 145989
rect 33567 145961 33601 145989
rect 33629 145961 33663 145989
rect 33691 145961 47619 145989
rect 47647 145961 47681 145989
rect 47709 145961 48837 145989
rect 48865 145961 48899 145989
rect 48927 145961 48961 145989
rect 48989 145961 49023 145989
rect 49051 145961 62979 145989
rect 63007 145961 63041 145989
rect 63069 145961 64197 145989
rect 64225 145961 64259 145989
rect 64287 145961 64321 145989
rect 64349 145961 64383 145989
rect 64411 145961 78339 145989
rect 78367 145961 78401 145989
rect 78429 145961 79557 145989
rect 79585 145961 79619 145989
rect 79647 145961 79681 145989
rect 79709 145961 79743 145989
rect 79771 145961 93699 145989
rect 93727 145961 93761 145989
rect 93789 145961 94917 145989
rect 94945 145961 94979 145989
rect 95007 145961 95041 145989
rect 95069 145961 95103 145989
rect 95131 145961 109059 145989
rect 109087 145961 109121 145989
rect 109149 145961 124419 145989
rect 124447 145961 124481 145989
rect 124509 145961 139779 145989
rect 139807 145961 139841 145989
rect 139869 145961 155139 145989
rect 155167 145961 155201 145989
rect 155229 145961 170499 145989
rect 170527 145961 170561 145989
rect 170589 145961 185859 145989
rect 185887 145961 185921 145989
rect 185949 145961 201219 145989
rect 201247 145961 201281 145989
rect 201309 145961 216579 145989
rect 216607 145961 216641 145989
rect 216669 145961 217797 145989
rect 217825 145961 217859 145989
rect 217887 145961 217921 145989
rect 217949 145961 217983 145989
rect 218011 145961 231939 145989
rect 231967 145961 232001 145989
rect 232029 145961 233157 145989
rect 233185 145961 233219 145989
rect 233247 145961 233281 145989
rect 233309 145961 233343 145989
rect 233371 145961 247299 145989
rect 247327 145961 247361 145989
rect 247389 145961 248517 145989
rect 248545 145961 248579 145989
rect 248607 145961 248641 145989
rect 248669 145961 248703 145989
rect 248731 145961 262659 145989
rect 262687 145961 262721 145989
rect 262749 145961 263877 145989
rect 263905 145961 263939 145989
rect 263967 145961 264001 145989
rect 264029 145961 264063 145989
rect 264091 145961 279237 145989
rect 279265 145961 279299 145989
rect 279327 145961 279361 145989
rect 279389 145961 279423 145989
rect 279451 145961 294597 145989
rect 294625 145961 294659 145989
rect 294687 145961 294721 145989
rect 294749 145961 294783 145989
rect 294811 145961 298248 145989
rect 298276 145961 298310 145989
rect 298338 145961 298372 145989
rect 298400 145961 298434 145989
rect 298462 145961 298990 145989
rect -958 145913 298990 145961
rect -958 140175 298990 140223
rect -958 140147 -910 140175
rect -882 140147 -848 140175
rect -820 140147 -786 140175
rect -758 140147 -724 140175
rect -696 140147 4617 140175
rect 4645 140147 4679 140175
rect 4707 140147 4741 140175
rect 4769 140147 4803 140175
rect 4831 140147 19977 140175
rect 20005 140147 20039 140175
rect 20067 140147 20101 140175
rect 20129 140147 20163 140175
rect 20191 140147 35337 140175
rect 35365 140147 35399 140175
rect 35427 140147 35461 140175
rect 35489 140147 35523 140175
rect 35551 140147 39939 140175
rect 39967 140147 40001 140175
rect 40029 140147 50697 140175
rect 50725 140147 50759 140175
rect 50787 140147 50821 140175
rect 50849 140147 50883 140175
rect 50911 140147 55299 140175
rect 55327 140147 55361 140175
rect 55389 140147 66057 140175
rect 66085 140147 66119 140175
rect 66147 140147 66181 140175
rect 66209 140147 66243 140175
rect 66271 140147 70659 140175
rect 70687 140147 70721 140175
rect 70749 140147 81417 140175
rect 81445 140147 81479 140175
rect 81507 140147 81541 140175
rect 81569 140147 81603 140175
rect 81631 140147 86019 140175
rect 86047 140147 86081 140175
rect 86109 140147 96777 140175
rect 96805 140147 96839 140175
rect 96867 140147 96901 140175
rect 96929 140147 96963 140175
rect 96991 140147 101379 140175
rect 101407 140147 101441 140175
rect 101469 140147 116739 140175
rect 116767 140147 116801 140175
rect 116829 140147 132099 140175
rect 132127 140147 132161 140175
rect 132189 140147 147459 140175
rect 147487 140147 147521 140175
rect 147549 140147 162819 140175
rect 162847 140147 162881 140175
rect 162909 140147 178179 140175
rect 178207 140147 178241 140175
rect 178269 140147 193539 140175
rect 193567 140147 193601 140175
rect 193629 140147 204297 140175
rect 204325 140147 204359 140175
rect 204387 140147 204421 140175
rect 204449 140147 204483 140175
rect 204511 140147 208899 140175
rect 208927 140147 208961 140175
rect 208989 140147 219657 140175
rect 219685 140147 219719 140175
rect 219747 140147 219781 140175
rect 219809 140147 219843 140175
rect 219871 140147 224259 140175
rect 224287 140147 224321 140175
rect 224349 140147 235017 140175
rect 235045 140147 235079 140175
rect 235107 140147 235141 140175
rect 235169 140147 235203 140175
rect 235231 140147 239619 140175
rect 239647 140147 239681 140175
rect 239709 140147 250377 140175
rect 250405 140147 250439 140175
rect 250467 140147 250501 140175
rect 250529 140147 250563 140175
rect 250591 140147 254979 140175
rect 255007 140147 255041 140175
rect 255069 140147 265737 140175
rect 265765 140147 265799 140175
rect 265827 140147 265861 140175
rect 265889 140147 265923 140175
rect 265951 140147 281097 140175
rect 281125 140147 281159 140175
rect 281187 140147 281221 140175
rect 281249 140147 281283 140175
rect 281311 140147 296457 140175
rect 296485 140147 296519 140175
rect 296547 140147 296581 140175
rect 296609 140147 296643 140175
rect 296671 140147 298728 140175
rect 298756 140147 298790 140175
rect 298818 140147 298852 140175
rect 298880 140147 298914 140175
rect 298942 140147 298990 140175
rect -958 140113 298990 140147
rect -958 140085 -910 140113
rect -882 140085 -848 140113
rect -820 140085 -786 140113
rect -758 140085 -724 140113
rect -696 140085 4617 140113
rect 4645 140085 4679 140113
rect 4707 140085 4741 140113
rect 4769 140085 4803 140113
rect 4831 140085 19977 140113
rect 20005 140085 20039 140113
rect 20067 140085 20101 140113
rect 20129 140085 20163 140113
rect 20191 140085 35337 140113
rect 35365 140085 35399 140113
rect 35427 140085 35461 140113
rect 35489 140085 35523 140113
rect 35551 140085 39939 140113
rect 39967 140085 40001 140113
rect 40029 140085 50697 140113
rect 50725 140085 50759 140113
rect 50787 140085 50821 140113
rect 50849 140085 50883 140113
rect 50911 140085 55299 140113
rect 55327 140085 55361 140113
rect 55389 140085 66057 140113
rect 66085 140085 66119 140113
rect 66147 140085 66181 140113
rect 66209 140085 66243 140113
rect 66271 140085 70659 140113
rect 70687 140085 70721 140113
rect 70749 140085 81417 140113
rect 81445 140085 81479 140113
rect 81507 140085 81541 140113
rect 81569 140085 81603 140113
rect 81631 140085 86019 140113
rect 86047 140085 86081 140113
rect 86109 140085 96777 140113
rect 96805 140085 96839 140113
rect 96867 140085 96901 140113
rect 96929 140085 96963 140113
rect 96991 140085 101379 140113
rect 101407 140085 101441 140113
rect 101469 140085 116739 140113
rect 116767 140085 116801 140113
rect 116829 140085 132099 140113
rect 132127 140085 132161 140113
rect 132189 140085 147459 140113
rect 147487 140085 147521 140113
rect 147549 140085 162819 140113
rect 162847 140085 162881 140113
rect 162909 140085 178179 140113
rect 178207 140085 178241 140113
rect 178269 140085 193539 140113
rect 193567 140085 193601 140113
rect 193629 140085 204297 140113
rect 204325 140085 204359 140113
rect 204387 140085 204421 140113
rect 204449 140085 204483 140113
rect 204511 140085 208899 140113
rect 208927 140085 208961 140113
rect 208989 140085 219657 140113
rect 219685 140085 219719 140113
rect 219747 140085 219781 140113
rect 219809 140085 219843 140113
rect 219871 140085 224259 140113
rect 224287 140085 224321 140113
rect 224349 140085 235017 140113
rect 235045 140085 235079 140113
rect 235107 140085 235141 140113
rect 235169 140085 235203 140113
rect 235231 140085 239619 140113
rect 239647 140085 239681 140113
rect 239709 140085 250377 140113
rect 250405 140085 250439 140113
rect 250467 140085 250501 140113
rect 250529 140085 250563 140113
rect 250591 140085 254979 140113
rect 255007 140085 255041 140113
rect 255069 140085 265737 140113
rect 265765 140085 265799 140113
rect 265827 140085 265861 140113
rect 265889 140085 265923 140113
rect 265951 140085 281097 140113
rect 281125 140085 281159 140113
rect 281187 140085 281221 140113
rect 281249 140085 281283 140113
rect 281311 140085 296457 140113
rect 296485 140085 296519 140113
rect 296547 140085 296581 140113
rect 296609 140085 296643 140113
rect 296671 140085 298728 140113
rect 298756 140085 298790 140113
rect 298818 140085 298852 140113
rect 298880 140085 298914 140113
rect 298942 140085 298990 140113
rect -958 140051 298990 140085
rect -958 140023 -910 140051
rect -882 140023 -848 140051
rect -820 140023 -786 140051
rect -758 140023 -724 140051
rect -696 140023 4617 140051
rect 4645 140023 4679 140051
rect 4707 140023 4741 140051
rect 4769 140023 4803 140051
rect 4831 140023 19977 140051
rect 20005 140023 20039 140051
rect 20067 140023 20101 140051
rect 20129 140023 20163 140051
rect 20191 140023 35337 140051
rect 35365 140023 35399 140051
rect 35427 140023 35461 140051
rect 35489 140023 35523 140051
rect 35551 140023 39939 140051
rect 39967 140023 40001 140051
rect 40029 140023 50697 140051
rect 50725 140023 50759 140051
rect 50787 140023 50821 140051
rect 50849 140023 50883 140051
rect 50911 140023 55299 140051
rect 55327 140023 55361 140051
rect 55389 140023 66057 140051
rect 66085 140023 66119 140051
rect 66147 140023 66181 140051
rect 66209 140023 66243 140051
rect 66271 140023 70659 140051
rect 70687 140023 70721 140051
rect 70749 140023 81417 140051
rect 81445 140023 81479 140051
rect 81507 140023 81541 140051
rect 81569 140023 81603 140051
rect 81631 140023 86019 140051
rect 86047 140023 86081 140051
rect 86109 140023 96777 140051
rect 96805 140023 96839 140051
rect 96867 140023 96901 140051
rect 96929 140023 96963 140051
rect 96991 140023 101379 140051
rect 101407 140023 101441 140051
rect 101469 140023 116739 140051
rect 116767 140023 116801 140051
rect 116829 140023 132099 140051
rect 132127 140023 132161 140051
rect 132189 140023 147459 140051
rect 147487 140023 147521 140051
rect 147549 140023 162819 140051
rect 162847 140023 162881 140051
rect 162909 140023 178179 140051
rect 178207 140023 178241 140051
rect 178269 140023 193539 140051
rect 193567 140023 193601 140051
rect 193629 140023 204297 140051
rect 204325 140023 204359 140051
rect 204387 140023 204421 140051
rect 204449 140023 204483 140051
rect 204511 140023 208899 140051
rect 208927 140023 208961 140051
rect 208989 140023 219657 140051
rect 219685 140023 219719 140051
rect 219747 140023 219781 140051
rect 219809 140023 219843 140051
rect 219871 140023 224259 140051
rect 224287 140023 224321 140051
rect 224349 140023 235017 140051
rect 235045 140023 235079 140051
rect 235107 140023 235141 140051
rect 235169 140023 235203 140051
rect 235231 140023 239619 140051
rect 239647 140023 239681 140051
rect 239709 140023 250377 140051
rect 250405 140023 250439 140051
rect 250467 140023 250501 140051
rect 250529 140023 250563 140051
rect 250591 140023 254979 140051
rect 255007 140023 255041 140051
rect 255069 140023 265737 140051
rect 265765 140023 265799 140051
rect 265827 140023 265861 140051
rect 265889 140023 265923 140051
rect 265951 140023 281097 140051
rect 281125 140023 281159 140051
rect 281187 140023 281221 140051
rect 281249 140023 281283 140051
rect 281311 140023 296457 140051
rect 296485 140023 296519 140051
rect 296547 140023 296581 140051
rect 296609 140023 296643 140051
rect 296671 140023 298728 140051
rect 298756 140023 298790 140051
rect 298818 140023 298852 140051
rect 298880 140023 298914 140051
rect 298942 140023 298990 140051
rect -958 139989 298990 140023
rect -958 139961 -910 139989
rect -882 139961 -848 139989
rect -820 139961 -786 139989
rect -758 139961 -724 139989
rect -696 139961 4617 139989
rect 4645 139961 4679 139989
rect 4707 139961 4741 139989
rect 4769 139961 4803 139989
rect 4831 139961 19977 139989
rect 20005 139961 20039 139989
rect 20067 139961 20101 139989
rect 20129 139961 20163 139989
rect 20191 139961 35337 139989
rect 35365 139961 35399 139989
rect 35427 139961 35461 139989
rect 35489 139961 35523 139989
rect 35551 139961 39939 139989
rect 39967 139961 40001 139989
rect 40029 139961 50697 139989
rect 50725 139961 50759 139989
rect 50787 139961 50821 139989
rect 50849 139961 50883 139989
rect 50911 139961 55299 139989
rect 55327 139961 55361 139989
rect 55389 139961 66057 139989
rect 66085 139961 66119 139989
rect 66147 139961 66181 139989
rect 66209 139961 66243 139989
rect 66271 139961 70659 139989
rect 70687 139961 70721 139989
rect 70749 139961 81417 139989
rect 81445 139961 81479 139989
rect 81507 139961 81541 139989
rect 81569 139961 81603 139989
rect 81631 139961 86019 139989
rect 86047 139961 86081 139989
rect 86109 139961 96777 139989
rect 96805 139961 96839 139989
rect 96867 139961 96901 139989
rect 96929 139961 96963 139989
rect 96991 139961 101379 139989
rect 101407 139961 101441 139989
rect 101469 139961 116739 139989
rect 116767 139961 116801 139989
rect 116829 139961 132099 139989
rect 132127 139961 132161 139989
rect 132189 139961 147459 139989
rect 147487 139961 147521 139989
rect 147549 139961 162819 139989
rect 162847 139961 162881 139989
rect 162909 139961 178179 139989
rect 178207 139961 178241 139989
rect 178269 139961 193539 139989
rect 193567 139961 193601 139989
rect 193629 139961 204297 139989
rect 204325 139961 204359 139989
rect 204387 139961 204421 139989
rect 204449 139961 204483 139989
rect 204511 139961 208899 139989
rect 208927 139961 208961 139989
rect 208989 139961 219657 139989
rect 219685 139961 219719 139989
rect 219747 139961 219781 139989
rect 219809 139961 219843 139989
rect 219871 139961 224259 139989
rect 224287 139961 224321 139989
rect 224349 139961 235017 139989
rect 235045 139961 235079 139989
rect 235107 139961 235141 139989
rect 235169 139961 235203 139989
rect 235231 139961 239619 139989
rect 239647 139961 239681 139989
rect 239709 139961 250377 139989
rect 250405 139961 250439 139989
rect 250467 139961 250501 139989
rect 250529 139961 250563 139989
rect 250591 139961 254979 139989
rect 255007 139961 255041 139989
rect 255069 139961 265737 139989
rect 265765 139961 265799 139989
rect 265827 139961 265861 139989
rect 265889 139961 265923 139989
rect 265951 139961 281097 139989
rect 281125 139961 281159 139989
rect 281187 139961 281221 139989
rect 281249 139961 281283 139989
rect 281311 139961 296457 139989
rect 296485 139961 296519 139989
rect 296547 139961 296581 139989
rect 296609 139961 296643 139989
rect 296671 139961 298728 139989
rect 298756 139961 298790 139989
rect 298818 139961 298852 139989
rect 298880 139961 298914 139989
rect 298942 139961 298990 139989
rect -958 139913 298990 139961
rect -958 137175 298990 137223
rect -958 137147 -430 137175
rect -402 137147 -368 137175
rect -340 137147 -306 137175
rect -278 137147 -244 137175
rect -216 137147 2757 137175
rect 2785 137147 2819 137175
rect 2847 137147 2881 137175
rect 2909 137147 2943 137175
rect 2971 137147 18117 137175
rect 18145 137147 18179 137175
rect 18207 137147 18241 137175
rect 18269 137147 18303 137175
rect 18331 137147 32259 137175
rect 32287 137147 32321 137175
rect 32349 137147 33477 137175
rect 33505 137147 33539 137175
rect 33567 137147 33601 137175
rect 33629 137147 33663 137175
rect 33691 137147 47619 137175
rect 47647 137147 47681 137175
rect 47709 137147 48837 137175
rect 48865 137147 48899 137175
rect 48927 137147 48961 137175
rect 48989 137147 49023 137175
rect 49051 137147 62979 137175
rect 63007 137147 63041 137175
rect 63069 137147 64197 137175
rect 64225 137147 64259 137175
rect 64287 137147 64321 137175
rect 64349 137147 64383 137175
rect 64411 137147 78339 137175
rect 78367 137147 78401 137175
rect 78429 137147 79557 137175
rect 79585 137147 79619 137175
rect 79647 137147 79681 137175
rect 79709 137147 79743 137175
rect 79771 137147 93699 137175
rect 93727 137147 93761 137175
rect 93789 137147 94917 137175
rect 94945 137147 94979 137175
rect 95007 137147 95041 137175
rect 95069 137147 95103 137175
rect 95131 137147 109059 137175
rect 109087 137147 109121 137175
rect 109149 137147 124419 137175
rect 124447 137147 124481 137175
rect 124509 137147 139779 137175
rect 139807 137147 139841 137175
rect 139869 137147 155139 137175
rect 155167 137147 155201 137175
rect 155229 137147 170499 137175
rect 170527 137147 170561 137175
rect 170589 137147 185859 137175
rect 185887 137147 185921 137175
rect 185949 137147 201219 137175
rect 201247 137147 201281 137175
rect 201309 137147 216579 137175
rect 216607 137147 216641 137175
rect 216669 137147 217797 137175
rect 217825 137147 217859 137175
rect 217887 137147 217921 137175
rect 217949 137147 217983 137175
rect 218011 137147 231939 137175
rect 231967 137147 232001 137175
rect 232029 137147 233157 137175
rect 233185 137147 233219 137175
rect 233247 137147 233281 137175
rect 233309 137147 233343 137175
rect 233371 137147 247299 137175
rect 247327 137147 247361 137175
rect 247389 137147 248517 137175
rect 248545 137147 248579 137175
rect 248607 137147 248641 137175
rect 248669 137147 248703 137175
rect 248731 137147 262659 137175
rect 262687 137147 262721 137175
rect 262749 137147 263877 137175
rect 263905 137147 263939 137175
rect 263967 137147 264001 137175
rect 264029 137147 264063 137175
rect 264091 137147 279237 137175
rect 279265 137147 279299 137175
rect 279327 137147 279361 137175
rect 279389 137147 279423 137175
rect 279451 137147 294597 137175
rect 294625 137147 294659 137175
rect 294687 137147 294721 137175
rect 294749 137147 294783 137175
rect 294811 137147 298248 137175
rect 298276 137147 298310 137175
rect 298338 137147 298372 137175
rect 298400 137147 298434 137175
rect 298462 137147 298990 137175
rect -958 137113 298990 137147
rect -958 137085 -430 137113
rect -402 137085 -368 137113
rect -340 137085 -306 137113
rect -278 137085 -244 137113
rect -216 137085 2757 137113
rect 2785 137085 2819 137113
rect 2847 137085 2881 137113
rect 2909 137085 2943 137113
rect 2971 137085 18117 137113
rect 18145 137085 18179 137113
rect 18207 137085 18241 137113
rect 18269 137085 18303 137113
rect 18331 137085 32259 137113
rect 32287 137085 32321 137113
rect 32349 137085 33477 137113
rect 33505 137085 33539 137113
rect 33567 137085 33601 137113
rect 33629 137085 33663 137113
rect 33691 137085 47619 137113
rect 47647 137085 47681 137113
rect 47709 137085 48837 137113
rect 48865 137085 48899 137113
rect 48927 137085 48961 137113
rect 48989 137085 49023 137113
rect 49051 137085 62979 137113
rect 63007 137085 63041 137113
rect 63069 137085 64197 137113
rect 64225 137085 64259 137113
rect 64287 137085 64321 137113
rect 64349 137085 64383 137113
rect 64411 137085 78339 137113
rect 78367 137085 78401 137113
rect 78429 137085 79557 137113
rect 79585 137085 79619 137113
rect 79647 137085 79681 137113
rect 79709 137085 79743 137113
rect 79771 137085 93699 137113
rect 93727 137085 93761 137113
rect 93789 137085 94917 137113
rect 94945 137085 94979 137113
rect 95007 137085 95041 137113
rect 95069 137085 95103 137113
rect 95131 137085 109059 137113
rect 109087 137085 109121 137113
rect 109149 137085 124419 137113
rect 124447 137085 124481 137113
rect 124509 137085 139779 137113
rect 139807 137085 139841 137113
rect 139869 137085 155139 137113
rect 155167 137085 155201 137113
rect 155229 137085 170499 137113
rect 170527 137085 170561 137113
rect 170589 137085 185859 137113
rect 185887 137085 185921 137113
rect 185949 137085 201219 137113
rect 201247 137085 201281 137113
rect 201309 137085 216579 137113
rect 216607 137085 216641 137113
rect 216669 137085 217797 137113
rect 217825 137085 217859 137113
rect 217887 137085 217921 137113
rect 217949 137085 217983 137113
rect 218011 137085 231939 137113
rect 231967 137085 232001 137113
rect 232029 137085 233157 137113
rect 233185 137085 233219 137113
rect 233247 137085 233281 137113
rect 233309 137085 233343 137113
rect 233371 137085 247299 137113
rect 247327 137085 247361 137113
rect 247389 137085 248517 137113
rect 248545 137085 248579 137113
rect 248607 137085 248641 137113
rect 248669 137085 248703 137113
rect 248731 137085 262659 137113
rect 262687 137085 262721 137113
rect 262749 137085 263877 137113
rect 263905 137085 263939 137113
rect 263967 137085 264001 137113
rect 264029 137085 264063 137113
rect 264091 137085 279237 137113
rect 279265 137085 279299 137113
rect 279327 137085 279361 137113
rect 279389 137085 279423 137113
rect 279451 137085 294597 137113
rect 294625 137085 294659 137113
rect 294687 137085 294721 137113
rect 294749 137085 294783 137113
rect 294811 137085 298248 137113
rect 298276 137085 298310 137113
rect 298338 137085 298372 137113
rect 298400 137085 298434 137113
rect 298462 137085 298990 137113
rect -958 137051 298990 137085
rect -958 137023 -430 137051
rect -402 137023 -368 137051
rect -340 137023 -306 137051
rect -278 137023 -244 137051
rect -216 137023 2757 137051
rect 2785 137023 2819 137051
rect 2847 137023 2881 137051
rect 2909 137023 2943 137051
rect 2971 137023 18117 137051
rect 18145 137023 18179 137051
rect 18207 137023 18241 137051
rect 18269 137023 18303 137051
rect 18331 137023 32259 137051
rect 32287 137023 32321 137051
rect 32349 137023 33477 137051
rect 33505 137023 33539 137051
rect 33567 137023 33601 137051
rect 33629 137023 33663 137051
rect 33691 137023 47619 137051
rect 47647 137023 47681 137051
rect 47709 137023 48837 137051
rect 48865 137023 48899 137051
rect 48927 137023 48961 137051
rect 48989 137023 49023 137051
rect 49051 137023 62979 137051
rect 63007 137023 63041 137051
rect 63069 137023 64197 137051
rect 64225 137023 64259 137051
rect 64287 137023 64321 137051
rect 64349 137023 64383 137051
rect 64411 137023 78339 137051
rect 78367 137023 78401 137051
rect 78429 137023 79557 137051
rect 79585 137023 79619 137051
rect 79647 137023 79681 137051
rect 79709 137023 79743 137051
rect 79771 137023 93699 137051
rect 93727 137023 93761 137051
rect 93789 137023 94917 137051
rect 94945 137023 94979 137051
rect 95007 137023 95041 137051
rect 95069 137023 95103 137051
rect 95131 137023 109059 137051
rect 109087 137023 109121 137051
rect 109149 137023 124419 137051
rect 124447 137023 124481 137051
rect 124509 137023 139779 137051
rect 139807 137023 139841 137051
rect 139869 137023 155139 137051
rect 155167 137023 155201 137051
rect 155229 137023 170499 137051
rect 170527 137023 170561 137051
rect 170589 137023 185859 137051
rect 185887 137023 185921 137051
rect 185949 137023 201219 137051
rect 201247 137023 201281 137051
rect 201309 137023 216579 137051
rect 216607 137023 216641 137051
rect 216669 137023 217797 137051
rect 217825 137023 217859 137051
rect 217887 137023 217921 137051
rect 217949 137023 217983 137051
rect 218011 137023 231939 137051
rect 231967 137023 232001 137051
rect 232029 137023 233157 137051
rect 233185 137023 233219 137051
rect 233247 137023 233281 137051
rect 233309 137023 233343 137051
rect 233371 137023 247299 137051
rect 247327 137023 247361 137051
rect 247389 137023 248517 137051
rect 248545 137023 248579 137051
rect 248607 137023 248641 137051
rect 248669 137023 248703 137051
rect 248731 137023 262659 137051
rect 262687 137023 262721 137051
rect 262749 137023 263877 137051
rect 263905 137023 263939 137051
rect 263967 137023 264001 137051
rect 264029 137023 264063 137051
rect 264091 137023 279237 137051
rect 279265 137023 279299 137051
rect 279327 137023 279361 137051
rect 279389 137023 279423 137051
rect 279451 137023 294597 137051
rect 294625 137023 294659 137051
rect 294687 137023 294721 137051
rect 294749 137023 294783 137051
rect 294811 137023 298248 137051
rect 298276 137023 298310 137051
rect 298338 137023 298372 137051
rect 298400 137023 298434 137051
rect 298462 137023 298990 137051
rect -958 136989 298990 137023
rect -958 136961 -430 136989
rect -402 136961 -368 136989
rect -340 136961 -306 136989
rect -278 136961 -244 136989
rect -216 136961 2757 136989
rect 2785 136961 2819 136989
rect 2847 136961 2881 136989
rect 2909 136961 2943 136989
rect 2971 136961 18117 136989
rect 18145 136961 18179 136989
rect 18207 136961 18241 136989
rect 18269 136961 18303 136989
rect 18331 136961 32259 136989
rect 32287 136961 32321 136989
rect 32349 136961 33477 136989
rect 33505 136961 33539 136989
rect 33567 136961 33601 136989
rect 33629 136961 33663 136989
rect 33691 136961 47619 136989
rect 47647 136961 47681 136989
rect 47709 136961 48837 136989
rect 48865 136961 48899 136989
rect 48927 136961 48961 136989
rect 48989 136961 49023 136989
rect 49051 136961 62979 136989
rect 63007 136961 63041 136989
rect 63069 136961 64197 136989
rect 64225 136961 64259 136989
rect 64287 136961 64321 136989
rect 64349 136961 64383 136989
rect 64411 136961 78339 136989
rect 78367 136961 78401 136989
rect 78429 136961 79557 136989
rect 79585 136961 79619 136989
rect 79647 136961 79681 136989
rect 79709 136961 79743 136989
rect 79771 136961 93699 136989
rect 93727 136961 93761 136989
rect 93789 136961 94917 136989
rect 94945 136961 94979 136989
rect 95007 136961 95041 136989
rect 95069 136961 95103 136989
rect 95131 136961 109059 136989
rect 109087 136961 109121 136989
rect 109149 136961 124419 136989
rect 124447 136961 124481 136989
rect 124509 136961 139779 136989
rect 139807 136961 139841 136989
rect 139869 136961 155139 136989
rect 155167 136961 155201 136989
rect 155229 136961 170499 136989
rect 170527 136961 170561 136989
rect 170589 136961 185859 136989
rect 185887 136961 185921 136989
rect 185949 136961 201219 136989
rect 201247 136961 201281 136989
rect 201309 136961 216579 136989
rect 216607 136961 216641 136989
rect 216669 136961 217797 136989
rect 217825 136961 217859 136989
rect 217887 136961 217921 136989
rect 217949 136961 217983 136989
rect 218011 136961 231939 136989
rect 231967 136961 232001 136989
rect 232029 136961 233157 136989
rect 233185 136961 233219 136989
rect 233247 136961 233281 136989
rect 233309 136961 233343 136989
rect 233371 136961 247299 136989
rect 247327 136961 247361 136989
rect 247389 136961 248517 136989
rect 248545 136961 248579 136989
rect 248607 136961 248641 136989
rect 248669 136961 248703 136989
rect 248731 136961 262659 136989
rect 262687 136961 262721 136989
rect 262749 136961 263877 136989
rect 263905 136961 263939 136989
rect 263967 136961 264001 136989
rect 264029 136961 264063 136989
rect 264091 136961 279237 136989
rect 279265 136961 279299 136989
rect 279327 136961 279361 136989
rect 279389 136961 279423 136989
rect 279451 136961 294597 136989
rect 294625 136961 294659 136989
rect 294687 136961 294721 136989
rect 294749 136961 294783 136989
rect 294811 136961 298248 136989
rect 298276 136961 298310 136989
rect 298338 136961 298372 136989
rect 298400 136961 298434 136989
rect 298462 136961 298990 136989
rect -958 136913 298990 136961
rect -958 131175 298990 131223
rect -958 131147 -910 131175
rect -882 131147 -848 131175
rect -820 131147 -786 131175
rect -758 131147 -724 131175
rect -696 131147 4617 131175
rect 4645 131147 4679 131175
rect 4707 131147 4741 131175
rect 4769 131147 4803 131175
rect 4831 131147 19977 131175
rect 20005 131147 20039 131175
rect 20067 131147 20101 131175
rect 20129 131147 20163 131175
rect 20191 131147 35337 131175
rect 35365 131147 35399 131175
rect 35427 131147 35461 131175
rect 35489 131147 35523 131175
rect 35551 131147 50697 131175
rect 50725 131147 50759 131175
rect 50787 131147 50821 131175
rect 50849 131147 50883 131175
rect 50911 131147 66057 131175
rect 66085 131147 66119 131175
rect 66147 131147 66181 131175
rect 66209 131147 66243 131175
rect 66271 131147 81417 131175
rect 81445 131147 81479 131175
rect 81507 131147 81541 131175
rect 81569 131147 81603 131175
rect 81631 131147 96777 131175
rect 96805 131147 96839 131175
rect 96867 131147 96901 131175
rect 96929 131147 96963 131175
rect 96991 131147 204297 131175
rect 204325 131147 204359 131175
rect 204387 131147 204421 131175
rect 204449 131147 204483 131175
rect 204511 131147 219657 131175
rect 219685 131147 219719 131175
rect 219747 131147 219781 131175
rect 219809 131147 219843 131175
rect 219871 131147 235017 131175
rect 235045 131147 235079 131175
rect 235107 131147 235141 131175
rect 235169 131147 235203 131175
rect 235231 131147 250377 131175
rect 250405 131147 250439 131175
rect 250467 131147 250501 131175
rect 250529 131147 250563 131175
rect 250591 131147 265737 131175
rect 265765 131147 265799 131175
rect 265827 131147 265861 131175
rect 265889 131147 265923 131175
rect 265951 131147 281097 131175
rect 281125 131147 281159 131175
rect 281187 131147 281221 131175
rect 281249 131147 281283 131175
rect 281311 131147 296457 131175
rect 296485 131147 296519 131175
rect 296547 131147 296581 131175
rect 296609 131147 296643 131175
rect 296671 131147 298728 131175
rect 298756 131147 298790 131175
rect 298818 131147 298852 131175
rect 298880 131147 298914 131175
rect 298942 131147 298990 131175
rect -958 131113 298990 131147
rect -958 131085 -910 131113
rect -882 131085 -848 131113
rect -820 131085 -786 131113
rect -758 131085 -724 131113
rect -696 131085 4617 131113
rect 4645 131085 4679 131113
rect 4707 131085 4741 131113
rect 4769 131085 4803 131113
rect 4831 131085 19977 131113
rect 20005 131085 20039 131113
rect 20067 131085 20101 131113
rect 20129 131085 20163 131113
rect 20191 131085 35337 131113
rect 35365 131085 35399 131113
rect 35427 131085 35461 131113
rect 35489 131085 35523 131113
rect 35551 131085 50697 131113
rect 50725 131085 50759 131113
rect 50787 131085 50821 131113
rect 50849 131085 50883 131113
rect 50911 131085 66057 131113
rect 66085 131085 66119 131113
rect 66147 131085 66181 131113
rect 66209 131085 66243 131113
rect 66271 131085 81417 131113
rect 81445 131085 81479 131113
rect 81507 131085 81541 131113
rect 81569 131085 81603 131113
rect 81631 131085 96777 131113
rect 96805 131085 96839 131113
rect 96867 131085 96901 131113
rect 96929 131085 96963 131113
rect 96991 131085 204297 131113
rect 204325 131085 204359 131113
rect 204387 131085 204421 131113
rect 204449 131085 204483 131113
rect 204511 131085 219657 131113
rect 219685 131085 219719 131113
rect 219747 131085 219781 131113
rect 219809 131085 219843 131113
rect 219871 131085 235017 131113
rect 235045 131085 235079 131113
rect 235107 131085 235141 131113
rect 235169 131085 235203 131113
rect 235231 131085 250377 131113
rect 250405 131085 250439 131113
rect 250467 131085 250501 131113
rect 250529 131085 250563 131113
rect 250591 131085 265737 131113
rect 265765 131085 265799 131113
rect 265827 131085 265861 131113
rect 265889 131085 265923 131113
rect 265951 131085 281097 131113
rect 281125 131085 281159 131113
rect 281187 131085 281221 131113
rect 281249 131085 281283 131113
rect 281311 131085 296457 131113
rect 296485 131085 296519 131113
rect 296547 131085 296581 131113
rect 296609 131085 296643 131113
rect 296671 131085 298728 131113
rect 298756 131085 298790 131113
rect 298818 131085 298852 131113
rect 298880 131085 298914 131113
rect 298942 131085 298990 131113
rect -958 131051 298990 131085
rect -958 131023 -910 131051
rect -882 131023 -848 131051
rect -820 131023 -786 131051
rect -758 131023 -724 131051
rect -696 131023 4617 131051
rect 4645 131023 4679 131051
rect 4707 131023 4741 131051
rect 4769 131023 4803 131051
rect 4831 131023 19977 131051
rect 20005 131023 20039 131051
rect 20067 131023 20101 131051
rect 20129 131023 20163 131051
rect 20191 131023 35337 131051
rect 35365 131023 35399 131051
rect 35427 131023 35461 131051
rect 35489 131023 35523 131051
rect 35551 131023 50697 131051
rect 50725 131023 50759 131051
rect 50787 131023 50821 131051
rect 50849 131023 50883 131051
rect 50911 131023 66057 131051
rect 66085 131023 66119 131051
rect 66147 131023 66181 131051
rect 66209 131023 66243 131051
rect 66271 131023 81417 131051
rect 81445 131023 81479 131051
rect 81507 131023 81541 131051
rect 81569 131023 81603 131051
rect 81631 131023 96777 131051
rect 96805 131023 96839 131051
rect 96867 131023 96901 131051
rect 96929 131023 96963 131051
rect 96991 131023 204297 131051
rect 204325 131023 204359 131051
rect 204387 131023 204421 131051
rect 204449 131023 204483 131051
rect 204511 131023 219657 131051
rect 219685 131023 219719 131051
rect 219747 131023 219781 131051
rect 219809 131023 219843 131051
rect 219871 131023 235017 131051
rect 235045 131023 235079 131051
rect 235107 131023 235141 131051
rect 235169 131023 235203 131051
rect 235231 131023 250377 131051
rect 250405 131023 250439 131051
rect 250467 131023 250501 131051
rect 250529 131023 250563 131051
rect 250591 131023 265737 131051
rect 265765 131023 265799 131051
rect 265827 131023 265861 131051
rect 265889 131023 265923 131051
rect 265951 131023 281097 131051
rect 281125 131023 281159 131051
rect 281187 131023 281221 131051
rect 281249 131023 281283 131051
rect 281311 131023 296457 131051
rect 296485 131023 296519 131051
rect 296547 131023 296581 131051
rect 296609 131023 296643 131051
rect 296671 131023 298728 131051
rect 298756 131023 298790 131051
rect 298818 131023 298852 131051
rect 298880 131023 298914 131051
rect 298942 131023 298990 131051
rect -958 131014 298990 131023
rect -958 130989 112137 131014
rect -958 130961 -910 130989
rect -882 130961 -848 130989
rect -820 130961 -786 130989
rect -758 130961 -724 130989
rect -696 130961 4617 130989
rect 4645 130961 4679 130989
rect 4707 130961 4741 130989
rect 4769 130961 4803 130989
rect 4831 130961 19977 130989
rect 20005 130961 20039 130989
rect 20067 130961 20101 130989
rect 20129 130961 20163 130989
rect 20191 130961 35337 130989
rect 35365 130961 35399 130989
rect 35427 130961 35461 130989
rect 35489 130961 35523 130989
rect 35551 130961 50697 130989
rect 50725 130961 50759 130989
rect 50787 130961 50821 130989
rect 50849 130961 50883 130989
rect 50911 130961 66057 130989
rect 66085 130961 66119 130989
rect 66147 130961 66181 130989
rect 66209 130961 66243 130989
rect 66271 130961 81417 130989
rect 81445 130961 81479 130989
rect 81507 130961 81541 130989
rect 81569 130961 81603 130989
rect 81631 130961 96777 130989
rect 96805 130961 96839 130989
rect 96867 130961 96901 130989
rect 96929 130961 96963 130989
rect 96991 130986 112137 130989
rect 112165 130986 112199 131014
rect 112227 130986 112261 131014
rect 112289 130986 112323 131014
rect 112351 130986 127497 131014
rect 127525 130986 127559 131014
rect 127587 130986 127621 131014
rect 127649 130986 127683 131014
rect 127711 130986 142857 131014
rect 142885 130986 142919 131014
rect 142947 130986 142981 131014
rect 143009 130986 143043 131014
rect 143071 130986 158217 131014
rect 158245 130986 158279 131014
rect 158307 130986 158341 131014
rect 158369 130986 158403 131014
rect 158431 130986 173577 131014
rect 173605 130986 173639 131014
rect 173667 130986 173701 131014
rect 173729 130986 173763 131014
rect 173791 130986 188937 131014
rect 188965 130986 188999 131014
rect 189027 130986 189061 131014
rect 189089 130986 189123 131014
rect 189151 130989 298990 131014
rect 189151 130986 204297 130989
rect 96991 130961 204297 130986
rect 204325 130961 204359 130989
rect 204387 130961 204421 130989
rect 204449 130961 204483 130989
rect 204511 130961 219657 130989
rect 219685 130961 219719 130989
rect 219747 130961 219781 130989
rect 219809 130961 219843 130989
rect 219871 130961 235017 130989
rect 235045 130961 235079 130989
rect 235107 130961 235141 130989
rect 235169 130961 235203 130989
rect 235231 130961 250377 130989
rect 250405 130961 250439 130989
rect 250467 130961 250501 130989
rect 250529 130961 250563 130989
rect 250591 130961 265737 130989
rect 265765 130961 265799 130989
rect 265827 130961 265861 130989
rect 265889 130961 265923 130989
rect 265951 130961 281097 130989
rect 281125 130961 281159 130989
rect 281187 130961 281221 130989
rect 281249 130961 281283 130989
rect 281311 130961 296457 130989
rect 296485 130961 296519 130989
rect 296547 130961 296581 130989
rect 296609 130961 296643 130989
rect 296671 130961 298728 130989
rect 298756 130961 298790 130989
rect 298818 130961 298852 130989
rect 298880 130961 298914 130989
rect 298942 130961 298990 130989
rect -958 130952 298990 130961
rect -958 130924 112137 130952
rect 112165 130924 112199 130952
rect 112227 130924 112261 130952
rect 112289 130924 112323 130952
rect 112351 130924 127497 130952
rect 127525 130924 127559 130952
rect 127587 130924 127621 130952
rect 127649 130924 127683 130952
rect 127711 130924 142857 130952
rect 142885 130924 142919 130952
rect 142947 130924 142981 130952
rect 143009 130924 143043 130952
rect 143071 130924 158217 130952
rect 158245 130924 158279 130952
rect 158307 130924 158341 130952
rect 158369 130924 158403 130952
rect 158431 130924 173577 130952
rect 173605 130924 173639 130952
rect 173667 130924 173701 130952
rect 173729 130924 173763 130952
rect 173791 130924 188937 130952
rect 188965 130924 188999 130952
rect 189027 130924 189061 130952
rect 189089 130924 189123 130952
rect 189151 130924 298990 130952
rect -958 130913 298990 130924
rect -958 128175 298990 128223
rect -958 128147 -430 128175
rect -402 128147 -368 128175
rect -340 128147 -306 128175
rect -278 128147 -244 128175
rect -216 128147 2757 128175
rect 2785 128147 2819 128175
rect 2847 128147 2881 128175
rect 2909 128147 2943 128175
rect 2971 128147 18117 128175
rect 18145 128147 18179 128175
rect 18207 128147 18241 128175
rect 18269 128147 18303 128175
rect 18331 128147 33477 128175
rect 33505 128147 33539 128175
rect 33567 128147 33601 128175
rect 33629 128147 33663 128175
rect 33691 128147 48837 128175
rect 48865 128147 48899 128175
rect 48927 128147 48961 128175
rect 48989 128147 49023 128175
rect 49051 128147 64197 128175
rect 64225 128147 64259 128175
rect 64287 128147 64321 128175
rect 64349 128147 64383 128175
rect 64411 128147 79557 128175
rect 79585 128147 79619 128175
rect 79647 128147 79681 128175
rect 79709 128147 79743 128175
rect 79771 128147 94917 128175
rect 94945 128147 94979 128175
rect 95007 128147 95041 128175
rect 95069 128147 95103 128175
rect 95131 128147 125637 128175
rect 125665 128147 125699 128175
rect 125727 128147 125761 128175
rect 125789 128147 125823 128175
rect 125851 128147 140997 128175
rect 141025 128147 141059 128175
rect 141087 128147 141121 128175
rect 141149 128147 141183 128175
rect 141211 128147 156357 128175
rect 156385 128147 156419 128175
rect 156447 128147 156481 128175
rect 156509 128147 156543 128175
rect 156571 128147 217797 128175
rect 217825 128147 217859 128175
rect 217887 128147 217921 128175
rect 217949 128147 217983 128175
rect 218011 128147 233157 128175
rect 233185 128147 233219 128175
rect 233247 128147 233281 128175
rect 233309 128147 233343 128175
rect 233371 128147 248517 128175
rect 248545 128147 248579 128175
rect 248607 128147 248641 128175
rect 248669 128147 248703 128175
rect 248731 128147 263877 128175
rect 263905 128147 263939 128175
rect 263967 128147 264001 128175
rect 264029 128147 264063 128175
rect 264091 128147 279237 128175
rect 279265 128147 279299 128175
rect 279327 128147 279361 128175
rect 279389 128147 279423 128175
rect 279451 128147 294597 128175
rect 294625 128147 294659 128175
rect 294687 128147 294721 128175
rect 294749 128147 294783 128175
rect 294811 128147 298248 128175
rect 298276 128147 298310 128175
rect 298338 128147 298372 128175
rect 298400 128147 298434 128175
rect 298462 128147 298990 128175
rect -958 128113 298990 128147
rect -958 128085 -430 128113
rect -402 128085 -368 128113
rect -340 128085 -306 128113
rect -278 128085 -244 128113
rect -216 128085 2757 128113
rect 2785 128085 2819 128113
rect 2847 128085 2881 128113
rect 2909 128085 2943 128113
rect 2971 128085 18117 128113
rect 18145 128085 18179 128113
rect 18207 128085 18241 128113
rect 18269 128085 18303 128113
rect 18331 128085 33477 128113
rect 33505 128085 33539 128113
rect 33567 128085 33601 128113
rect 33629 128085 33663 128113
rect 33691 128085 48837 128113
rect 48865 128085 48899 128113
rect 48927 128085 48961 128113
rect 48989 128085 49023 128113
rect 49051 128085 64197 128113
rect 64225 128085 64259 128113
rect 64287 128085 64321 128113
rect 64349 128085 64383 128113
rect 64411 128085 79557 128113
rect 79585 128085 79619 128113
rect 79647 128085 79681 128113
rect 79709 128085 79743 128113
rect 79771 128085 94917 128113
rect 94945 128085 94979 128113
rect 95007 128085 95041 128113
rect 95069 128085 95103 128113
rect 95131 128085 125637 128113
rect 125665 128085 125699 128113
rect 125727 128085 125761 128113
rect 125789 128085 125823 128113
rect 125851 128085 140997 128113
rect 141025 128085 141059 128113
rect 141087 128085 141121 128113
rect 141149 128085 141183 128113
rect 141211 128085 156357 128113
rect 156385 128085 156419 128113
rect 156447 128085 156481 128113
rect 156509 128085 156543 128113
rect 156571 128085 217797 128113
rect 217825 128085 217859 128113
rect 217887 128085 217921 128113
rect 217949 128085 217983 128113
rect 218011 128085 233157 128113
rect 233185 128085 233219 128113
rect 233247 128085 233281 128113
rect 233309 128085 233343 128113
rect 233371 128085 248517 128113
rect 248545 128085 248579 128113
rect 248607 128085 248641 128113
rect 248669 128085 248703 128113
rect 248731 128085 263877 128113
rect 263905 128085 263939 128113
rect 263967 128085 264001 128113
rect 264029 128085 264063 128113
rect 264091 128085 279237 128113
rect 279265 128085 279299 128113
rect 279327 128085 279361 128113
rect 279389 128085 279423 128113
rect 279451 128085 294597 128113
rect 294625 128085 294659 128113
rect 294687 128085 294721 128113
rect 294749 128085 294783 128113
rect 294811 128085 298248 128113
rect 298276 128085 298310 128113
rect 298338 128085 298372 128113
rect 298400 128085 298434 128113
rect 298462 128085 298990 128113
rect -958 128051 298990 128085
rect -958 128023 -430 128051
rect -402 128023 -368 128051
rect -340 128023 -306 128051
rect -278 128023 -244 128051
rect -216 128023 2757 128051
rect 2785 128023 2819 128051
rect 2847 128023 2881 128051
rect 2909 128023 2943 128051
rect 2971 128023 18117 128051
rect 18145 128023 18179 128051
rect 18207 128023 18241 128051
rect 18269 128023 18303 128051
rect 18331 128023 33477 128051
rect 33505 128023 33539 128051
rect 33567 128023 33601 128051
rect 33629 128023 33663 128051
rect 33691 128023 48837 128051
rect 48865 128023 48899 128051
rect 48927 128023 48961 128051
rect 48989 128023 49023 128051
rect 49051 128023 64197 128051
rect 64225 128023 64259 128051
rect 64287 128023 64321 128051
rect 64349 128023 64383 128051
rect 64411 128023 79557 128051
rect 79585 128023 79619 128051
rect 79647 128023 79681 128051
rect 79709 128023 79743 128051
rect 79771 128023 94917 128051
rect 94945 128023 94979 128051
rect 95007 128023 95041 128051
rect 95069 128023 95103 128051
rect 95131 128023 125637 128051
rect 125665 128023 125699 128051
rect 125727 128023 125761 128051
rect 125789 128023 125823 128051
rect 125851 128023 140997 128051
rect 141025 128023 141059 128051
rect 141087 128023 141121 128051
rect 141149 128023 141183 128051
rect 141211 128023 156357 128051
rect 156385 128023 156419 128051
rect 156447 128023 156481 128051
rect 156509 128023 156543 128051
rect 156571 128023 217797 128051
rect 217825 128023 217859 128051
rect 217887 128023 217921 128051
rect 217949 128023 217983 128051
rect 218011 128023 233157 128051
rect 233185 128023 233219 128051
rect 233247 128023 233281 128051
rect 233309 128023 233343 128051
rect 233371 128023 248517 128051
rect 248545 128023 248579 128051
rect 248607 128023 248641 128051
rect 248669 128023 248703 128051
rect 248731 128023 263877 128051
rect 263905 128023 263939 128051
rect 263967 128023 264001 128051
rect 264029 128023 264063 128051
rect 264091 128023 279237 128051
rect 279265 128023 279299 128051
rect 279327 128023 279361 128051
rect 279389 128023 279423 128051
rect 279451 128023 294597 128051
rect 294625 128023 294659 128051
rect 294687 128023 294721 128051
rect 294749 128023 294783 128051
rect 294811 128023 298248 128051
rect 298276 128023 298310 128051
rect 298338 128023 298372 128051
rect 298400 128023 298434 128051
rect 298462 128023 298990 128051
rect -958 127989 298990 128023
rect -958 127961 -430 127989
rect -402 127961 -368 127989
rect -340 127961 -306 127989
rect -278 127961 -244 127989
rect -216 127961 2757 127989
rect 2785 127961 2819 127989
rect 2847 127961 2881 127989
rect 2909 127961 2943 127989
rect 2971 127961 18117 127989
rect 18145 127961 18179 127989
rect 18207 127961 18241 127989
rect 18269 127961 18303 127989
rect 18331 127961 33477 127989
rect 33505 127961 33539 127989
rect 33567 127961 33601 127989
rect 33629 127961 33663 127989
rect 33691 127961 48837 127989
rect 48865 127961 48899 127989
rect 48927 127961 48961 127989
rect 48989 127961 49023 127989
rect 49051 127961 64197 127989
rect 64225 127961 64259 127989
rect 64287 127961 64321 127989
rect 64349 127961 64383 127989
rect 64411 127961 79557 127989
rect 79585 127961 79619 127989
rect 79647 127961 79681 127989
rect 79709 127961 79743 127989
rect 79771 127961 94917 127989
rect 94945 127961 94979 127989
rect 95007 127961 95041 127989
rect 95069 127961 95103 127989
rect 95131 127961 125637 127989
rect 125665 127961 125699 127989
rect 125727 127961 125761 127989
rect 125789 127961 125823 127989
rect 125851 127961 140997 127989
rect 141025 127961 141059 127989
rect 141087 127961 141121 127989
rect 141149 127961 141183 127989
rect 141211 127961 156357 127989
rect 156385 127961 156419 127989
rect 156447 127961 156481 127989
rect 156509 127961 156543 127989
rect 156571 127961 217797 127989
rect 217825 127961 217859 127989
rect 217887 127961 217921 127989
rect 217949 127961 217983 127989
rect 218011 127961 233157 127989
rect 233185 127961 233219 127989
rect 233247 127961 233281 127989
rect 233309 127961 233343 127989
rect 233371 127961 248517 127989
rect 248545 127961 248579 127989
rect 248607 127961 248641 127989
rect 248669 127961 248703 127989
rect 248731 127961 263877 127989
rect 263905 127961 263939 127989
rect 263967 127961 264001 127989
rect 264029 127961 264063 127989
rect 264091 127961 279237 127989
rect 279265 127961 279299 127989
rect 279327 127961 279361 127989
rect 279389 127961 279423 127989
rect 279451 127961 294597 127989
rect 294625 127961 294659 127989
rect 294687 127961 294721 127989
rect 294749 127961 294783 127989
rect 294811 127961 298248 127989
rect 298276 127961 298310 127989
rect 298338 127961 298372 127989
rect 298400 127961 298434 127989
rect 298462 127961 298990 127989
rect -958 127913 298990 127961
rect -958 122175 298990 122223
rect -958 122147 -910 122175
rect -882 122147 -848 122175
rect -820 122147 -786 122175
rect -758 122147 -724 122175
rect -696 122147 4617 122175
rect 4645 122147 4679 122175
rect 4707 122147 4741 122175
rect 4769 122147 4803 122175
rect 4831 122147 19977 122175
rect 20005 122147 20039 122175
rect 20067 122147 20101 122175
rect 20129 122147 20163 122175
rect 20191 122147 35337 122175
rect 35365 122147 35399 122175
rect 35427 122147 35461 122175
rect 35489 122147 35523 122175
rect 35551 122147 50697 122175
rect 50725 122147 50759 122175
rect 50787 122147 50821 122175
rect 50849 122147 50883 122175
rect 50911 122147 66057 122175
rect 66085 122147 66119 122175
rect 66147 122147 66181 122175
rect 66209 122147 66243 122175
rect 66271 122147 81417 122175
rect 81445 122147 81479 122175
rect 81507 122147 81541 122175
rect 81569 122147 81603 122175
rect 81631 122147 96777 122175
rect 96805 122147 96839 122175
rect 96867 122147 96901 122175
rect 96929 122147 96963 122175
rect 96991 122147 109939 122175
rect 109967 122147 110001 122175
rect 110029 122147 112137 122175
rect 112165 122147 112199 122175
rect 112227 122147 112261 122175
rect 112289 122147 112323 122175
rect 112351 122147 125299 122175
rect 125327 122147 125361 122175
rect 125389 122147 127497 122175
rect 127525 122147 127559 122175
rect 127587 122147 127621 122175
rect 127649 122147 127683 122175
rect 127711 122147 142857 122175
rect 142885 122147 142919 122175
rect 142947 122147 142981 122175
rect 143009 122147 143043 122175
rect 143071 122147 158217 122175
rect 158245 122147 158279 122175
rect 158307 122147 158341 122175
rect 158369 122147 158403 122175
rect 158431 122147 169939 122175
rect 169967 122147 170001 122175
rect 170029 122147 185299 122175
rect 185327 122147 185361 122175
rect 185389 122147 200659 122175
rect 200687 122147 200721 122175
rect 200749 122147 216019 122175
rect 216047 122147 216081 122175
rect 216109 122147 231379 122175
rect 231407 122147 231441 122175
rect 231469 122147 246739 122175
rect 246767 122147 246801 122175
rect 246829 122147 262099 122175
rect 262127 122147 262161 122175
rect 262189 122147 281097 122175
rect 281125 122147 281159 122175
rect 281187 122147 281221 122175
rect 281249 122147 281283 122175
rect 281311 122147 296457 122175
rect 296485 122147 296519 122175
rect 296547 122147 296581 122175
rect 296609 122147 296643 122175
rect 296671 122147 298728 122175
rect 298756 122147 298790 122175
rect 298818 122147 298852 122175
rect 298880 122147 298914 122175
rect 298942 122147 298990 122175
rect -958 122113 298990 122147
rect -958 122085 -910 122113
rect -882 122085 -848 122113
rect -820 122085 -786 122113
rect -758 122085 -724 122113
rect -696 122085 4617 122113
rect 4645 122085 4679 122113
rect 4707 122085 4741 122113
rect 4769 122085 4803 122113
rect 4831 122085 19977 122113
rect 20005 122085 20039 122113
rect 20067 122085 20101 122113
rect 20129 122085 20163 122113
rect 20191 122085 35337 122113
rect 35365 122085 35399 122113
rect 35427 122085 35461 122113
rect 35489 122085 35523 122113
rect 35551 122085 50697 122113
rect 50725 122085 50759 122113
rect 50787 122085 50821 122113
rect 50849 122085 50883 122113
rect 50911 122085 66057 122113
rect 66085 122085 66119 122113
rect 66147 122085 66181 122113
rect 66209 122085 66243 122113
rect 66271 122085 81417 122113
rect 81445 122085 81479 122113
rect 81507 122085 81541 122113
rect 81569 122085 81603 122113
rect 81631 122085 96777 122113
rect 96805 122085 96839 122113
rect 96867 122085 96901 122113
rect 96929 122085 96963 122113
rect 96991 122085 109939 122113
rect 109967 122085 110001 122113
rect 110029 122085 112137 122113
rect 112165 122085 112199 122113
rect 112227 122085 112261 122113
rect 112289 122085 112323 122113
rect 112351 122085 125299 122113
rect 125327 122085 125361 122113
rect 125389 122085 127497 122113
rect 127525 122085 127559 122113
rect 127587 122085 127621 122113
rect 127649 122085 127683 122113
rect 127711 122085 142857 122113
rect 142885 122085 142919 122113
rect 142947 122085 142981 122113
rect 143009 122085 143043 122113
rect 143071 122085 158217 122113
rect 158245 122085 158279 122113
rect 158307 122085 158341 122113
rect 158369 122085 158403 122113
rect 158431 122085 169939 122113
rect 169967 122085 170001 122113
rect 170029 122085 185299 122113
rect 185327 122085 185361 122113
rect 185389 122085 200659 122113
rect 200687 122085 200721 122113
rect 200749 122085 216019 122113
rect 216047 122085 216081 122113
rect 216109 122085 231379 122113
rect 231407 122085 231441 122113
rect 231469 122085 246739 122113
rect 246767 122085 246801 122113
rect 246829 122085 262099 122113
rect 262127 122085 262161 122113
rect 262189 122085 281097 122113
rect 281125 122085 281159 122113
rect 281187 122085 281221 122113
rect 281249 122085 281283 122113
rect 281311 122085 296457 122113
rect 296485 122085 296519 122113
rect 296547 122085 296581 122113
rect 296609 122085 296643 122113
rect 296671 122085 298728 122113
rect 298756 122085 298790 122113
rect 298818 122085 298852 122113
rect 298880 122085 298914 122113
rect 298942 122085 298990 122113
rect -958 122051 298990 122085
rect -958 122023 -910 122051
rect -882 122023 -848 122051
rect -820 122023 -786 122051
rect -758 122023 -724 122051
rect -696 122023 4617 122051
rect 4645 122023 4679 122051
rect 4707 122023 4741 122051
rect 4769 122023 4803 122051
rect 4831 122023 19977 122051
rect 20005 122023 20039 122051
rect 20067 122023 20101 122051
rect 20129 122023 20163 122051
rect 20191 122023 35337 122051
rect 35365 122023 35399 122051
rect 35427 122023 35461 122051
rect 35489 122023 35523 122051
rect 35551 122023 50697 122051
rect 50725 122023 50759 122051
rect 50787 122023 50821 122051
rect 50849 122023 50883 122051
rect 50911 122023 66057 122051
rect 66085 122023 66119 122051
rect 66147 122023 66181 122051
rect 66209 122023 66243 122051
rect 66271 122023 81417 122051
rect 81445 122023 81479 122051
rect 81507 122023 81541 122051
rect 81569 122023 81603 122051
rect 81631 122023 96777 122051
rect 96805 122023 96839 122051
rect 96867 122023 96901 122051
rect 96929 122023 96963 122051
rect 96991 122023 109939 122051
rect 109967 122023 110001 122051
rect 110029 122023 112137 122051
rect 112165 122023 112199 122051
rect 112227 122023 112261 122051
rect 112289 122023 112323 122051
rect 112351 122023 125299 122051
rect 125327 122023 125361 122051
rect 125389 122023 127497 122051
rect 127525 122023 127559 122051
rect 127587 122023 127621 122051
rect 127649 122023 127683 122051
rect 127711 122023 142857 122051
rect 142885 122023 142919 122051
rect 142947 122023 142981 122051
rect 143009 122023 143043 122051
rect 143071 122023 158217 122051
rect 158245 122023 158279 122051
rect 158307 122023 158341 122051
rect 158369 122023 158403 122051
rect 158431 122023 169939 122051
rect 169967 122023 170001 122051
rect 170029 122023 185299 122051
rect 185327 122023 185361 122051
rect 185389 122023 200659 122051
rect 200687 122023 200721 122051
rect 200749 122023 216019 122051
rect 216047 122023 216081 122051
rect 216109 122023 231379 122051
rect 231407 122023 231441 122051
rect 231469 122023 246739 122051
rect 246767 122023 246801 122051
rect 246829 122023 262099 122051
rect 262127 122023 262161 122051
rect 262189 122023 281097 122051
rect 281125 122023 281159 122051
rect 281187 122023 281221 122051
rect 281249 122023 281283 122051
rect 281311 122023 296457 122051
rect 296485 122023 296519 122051
rect 296547 122023 296581 122051
rect 296609 122023 296643 122051
rect 296671 122023 298728 122051
rect 298756 122023 298790 122051
rect 298818 122023 298852 122051
rect 298880 122023 298914 122051
rect 298942 122023 298990 122051
rect -958 121989 298990 122023
rect -958 121961 -910 121989
rect -882 121961 -848 121989
rect -820 121961 -786 121989
rect -758 121961 -724 121989
rect -696 121961 4617 121989
rect 4645 121961 4679 121989
rect 4707 121961 4741 121989
rect 4769 121961 4803 121989
rect 4831 121961 19977 121989
rect 20005 121961 20039 121989
rect 20067 121961 20101 121989
rect 20129 121961 20163 121989
rect 20191 121961 35337 121989
rect 35365 121961 35399 121989
rect 35427 121961 35461 121989
rect 35489 121961 35523 121989
rect 35551 121961 50697 121989
rect 50725 121961 50759 121989
rect 50787 121961 50821 121989
rect 50849 121961 50883 121989
rect 50911 121961 66057 121989
rect 66085 121961 66119 121989
rect 66147 121961 66181 121989
rect 66209 121961 66243 121989
rect 66271 121961 81417 121989
rect 81445 121961 81479 121989
rect 81507 121961 81541 121989
rect 81569 121961 81603 121989
rect 81631 121961 96777 121989
rect 96805 121961 96839 121989
rect 96867 121961 96901 121989
rect 96929 121961 96963 121989
rect 96991 121961 109939 121989
rect 109967 121961 110001 121989
rect 110029 121961 112137 121989
rect 112165 121961 112199 121989
rect 112227 121961 112261 121989
rect 112289 121961 112323 121989
rect 112351 121961 125299 121989
rect 125327 121961 125361 121989
rect 125389 121961 127497 121989
rect 127525 121961 127559 121989
rect 127587 121961 127621 121989
rect 127649 121961 127683 121989
rect 127711 121961 142857 121989
rect 142885 121961 142919 121989
rect 142947 121961 142981 121989
rect 143009 121961 143043 121989
rect 143071 121961 158217 121989
rect 158245 121961 158279 121989
rect 158307 121961 158341 121989
rect 158369 121961 158403 121989
rect 158431 121961 169939 121989
rect 169967 121961 170001 121989
rect 170029 121961 185299 121989
rect 185327 121961 185361 121989
rect 185389 121961 200659 121989
rect 200687 121961 200721 121989
rect 200749 121961 216019 121989
rect 216047 121961 216081 121989
rect 216109 121961 231379 121989
rect 231407 121961 231441 121989
rect 231469 121961 246739 121989
rect 246767 121961 246801 121989
rect 246829 121961 262099 121989
rect 262127 121961 262161 121989
rect 262189 121961 281097 121989
rect 281125 121961 281159 121989
rect 281187 121961 281221 121989
rect 281249 121961 281283 121989
rect 281311 121961 296457 121989
rect 296485 121961 296519 121989
rect 296547 121961 296581 121989
rect 296609 121961 296643 121989
rect 296671 121961 298728 121989
rect 298756 121961 298790 121989
rect 298818 121961 298852 121989
rect 298880 121961 298914 121989
rect 298942 121961 298990 121989
rect -958 121913 298990 121961
rect -958 119175 298990 119223
rect -958 119147 -430 119175
rect -402 119147 -368 119175
rect -340 119147 -306 119175
rect -278 119147 -244 119175
rect -216 119147 2757 119175
rect 2785 119147 2819 119175
rect 2847 119147 2881 119175
rect 2909 119147 2943 119175
rect 2971 119147 18117 119175
rect 18145 119147 18179 119175
rect 18207 119147 18241 119175
rect 18269 119147 18303 119175
rect 18331 119147 33477 119175
rect 33505 119147 33539 119175
rect 33567 119147 33601 119175
rect 33629 119147 33663 119175
rect 33691 119147 48837 119175
rect 48865 119147 48899 119175
rect 48927 119147 48961 119175
rect 48989 119147 49023 119175
rect 49051 119147 64197 119175
rect 64225 119147 64259 119175
rect 64287 119147 64321 119175
rect 64349 119147 64383 119175
rect 64411 119147 79557 119175
rect 79585 119147 79619 119175
rect 79647 119147 79681 119175
rect 79709 119147 79743 119175
rect 79771 119147 94917 119175
rect 94945 119147 94979 119175
rect 95007 119147 95041 119175
rect 95069 119147 95103 119175
rect 95131 119147 102259 119175
rect 102287 119147 102321 119175
rect 102349 119147 117619 119175
rect 117647 119147 117681 119175
rect 117709 119147 125637 119175
rect 125665 119147 125699 119175
rect 125727 119147 125761 119175
rect 125789 119147 125823 119175
rect 125851 119147 140997 119175
rect 141025 119147 141059 119175
rect 141087 119147 141121 119175
rect 141149 119147 141183 119175
rect 141211 119147 156357 119175
rect 156385 119147 156419 119175
rect 156447 119147 156481 119175
rect 156509 119147 156543 119175
rect 156571 119147 162259 119175
rect 162287 119147 162321 119175
rect 162349 119147 177619 119175
rect 177647 119147 177681 119175
rect 177709 119147 192979 119175
rect 193007 119147 193041 119175
rect 193069 119147 208339 119175
rect 208367 119147 208401 119175
rect 208429 119147 223699 119175
rect 223727 119147 223761 119175
rect 223789 119147 239059 119175
rect 239087 119147 239121 119175
rect 239149 119147 254419 119175
rect 254447 119147 254481 119175
rect 254509 119147 269779 119175
rect 269807 119147 269841 119175
rect 269869 119147 279237 119175
rect 279265 119147 279299 119175
rect 279327 119147 279361 119175
rect 279389 119147 279423 119175
rect 279451 119147 294597 119175
rect 294625 119147 294659 119175
rect 294687 119147 294721 119175
rect 294749 119147 294783 119175
rect 294811 119147 298248 119175
rect 298276 119147 298310 119175
rect 298338 119147 298372 119175
rect 298400 119147 298434 119175
rect 298462 119147 298990 119175
rect -958 119113 298990 119147
rect -958 119085 -430 119113
rect -402 119085 -368 119113
rect -340 119085 -306 119113
rect -278 119085 -244 119113
rect -216 119085 2757 119113
rect 2785 119085 2819 119113
rect 2847 119085 2881 119113
rect 2909 119085 2943 119113
rect 2971 119085 18117 119113
rect 18145 119085 18179 119113
rect 18207 119085 18241 119113
rect 18269 119085 18303 119113
rect 18331 119085 33477 119113
rect 33505 119085 33539 119113
rect 33567 119085 33601 119113
rect 33629 119085 33663 119113
rect 33691 119085 48837 119113
rect 48865 119085 48899 119113
rect 48927 119085 48961 119113
rect 48989 119085 49023 119113
rect 49051 119085 64197 119113
rect 64225 119085 64259 119113
rect 64287 119085 64321 119113
rect 64349 119085 64383 119113
rect 64411 119085 79557 119113
rect 79585 119085 79619 119113
rect 79647 119085 79681 119113
rect 79709 119085 79743 119113
rect 79771 119085 94917 119113
rect 94945 119085 94979 119113
rect 95007 119085 95041 119113
rect 95069 119085 95103 119113
rect 95131 119085 102259 119113
rect 102287 119085 102321 119113
rect 102349 119085 117619 119113
rect 117647 119085 117681 119113
rect 117709 119085 125637 119113
rect 125665 119085 125699 119113
rect 125727 119085 125761 119113
rect 125789 119085 125823 119113
rect 125851 119085 140997 119113
rect 141025 119085 141059 119113
rect 141087 119085 141121 119113
rect 141149 119085 141183 119113
rect 141211 119085 156357 119113
rect 156385 119085 156419 119113
rect 156447 119085 156481 119113
rect 156509 119085 156543 119113
rect 156571 119085 162259 119113
rect 162287 119085 162321 119113
rect 162349 119085 177619 119113
rect 177647 119085 177681 119113
rect 177709 119085 192979 119113
rect 193007 119085 193041 119113
rect 193069 119085 208339 119113
rect 208367 119085 208401 119113
rect 208429 119085 223699 119113
rect 223727 119085 223761 119113
rect 223789 119085 239059 119113
rect 239087 119085 239121 119113
rect 239149 119085 254419 119113
rect 254447 119085 254481 119113
rect 254509 119085 269779 119113
rect 269807 119085 269841 119113
rect 269869 119085 279237 119113
rect 279265 119085 279299 119113
rect 279327 119085 279361 119113
rect 279389 119085 279423 119113
rect 279451 119085 294597 119113
rect 294625 119085 294659 119113
rect 294687 119085 294721 119113
rect 294749 119085 294783 119113
rect 294811 119085 298248 119113
rect 298276 119085 298310 119113
rect 298338 119085 298372 119113
rect 298400 119085 298434 119113
rect 298462 119085 298990 119113
rect -958 119051 298990 119085
rect -958 119023 -430 119051
rect -402 119023 -368 119051
rect -340 119023 -306 119051
rect -278 119023 -244 119051
rect -216 119023 2757 119051
rect 2785 119023 2819 119051
rect 2847 119023 2881 119051
rect 2909 119023 2943 119051
rect 2971 119023 18117 119051
rect 18145 119023 18179 119051
rect 18207 119023 18241 119051
rect 18269 119023 18303 119051
rect 18331 119023 33477 119051
rect 33505 119023 33539 119051
rect 33567 119023 33601 119051
rect 33629 119023 33663 119051
rect 33691 119023 48837 119051
rect 48865 119023 48899 119051
rect 48927 119023 48961 119051
rect 48989 119023 49023 119051
rect 49051 119023 64197 119051
rect 64225 119023 64259 119051
rect 64287 119023 64321 119051
rect 64349 119023 64383 119051
rect 64411 119023 79557 119051
rect 79585 119023 79619 119051
rect 79647 119023 79681 119051
rect 79709 119023 79743 119051
rect 79771 119023 94917 119051
rect 94945 119023 94979 119051
rect 95007 119023 95041 119051
rect 95069 119023 95103 119051
rect 95131 119023 102259 119051
rect 102287 119023 102321 119051
rect 102349 119023 117619 119051
rect 117647 119023 117681 119051
rect 117709 119023 125637 119051
rect 125665 119023 125699 119051
rect 125727 119023 125761 119051
rect 125789 119023 125823 119051
rect 125851 119023 140997 119051
rect 141025 119023 141059 119051
rect 141087 119023 141121 119051
rect 141149 119023 141183 119051
rect 141211 119023 156357 119051
rect 156385 119023 156419 119051
rect 156447 119023 156481 119051
rect 156509 119023 156543 119051
rect 156571 119023 162259 119051
rect 162287 119023 162321 119051
rect 162349 119023 177619 119051
rect 177647 119023 177681 119051
rect 177709 119023 192979 119051
rect 193007 119023 193041 119051
rect 193069 119023 208339 119051
rect 208367 119023 208401 119051
rect 208429 119023 223699 119051
rect 223727 119023 223761 119051
rect 223789 119023 239059 119051
rect 239087 119023 239121 119051
rect 239149 119023 254419 119051
rect 254447 119023 254481 119051
rect 254509 119023 269779 119051
rect 269807 119023 269841 119051
rect 269869 119023 279237 119051
rect 279265 119023 279299 119051
rect 279327 119023 279361 119051
rect 279389 119023 279423 119051
rect 279451 119023 294597 119051
rect 294625 119023 294659 119051
rect 294687 119023 294721 119051
rect 294749 119023 294783 119051
rect 294811 119023 298248 119051
rect 298276 119023 298310 119051
rect 298338 119023 298372 119051
rect 298400 119023 298434 119051
rect 298462 119023 298990 119051
rect -958 118989 298990 119023
rect -958 118961 -430 118989
rect -402 118961 -368 118989
rect -340 118961 -306 118989
rect -278 118961 -244 118989
rect -216 118961 2757 118989
rect 2785 118961 2819 118989
rect 2847 118961 2881 118989
rect 2909 118961 2943 118989
rect 2971 118961 18117 118989
rect 18145 118961 18179 118989
rect 18207 118961 18241 118989
rect 18269 118961 18303 118989
rect 18331 118961 33477 118989
rect 33505 118961 33539 118989
rect 33567 118961 33601 118989
rect 33629 118961 33663 118989
rect 33691 118961 48837 118989
rect 48865 118961 48899 118989
rect 48927 118961 48961 118989
rect 48989 118961 49023 118989
rect 49051 118961 64197 118989
rect 64225 118961 64259 118989
rect 64287 118961 64321 118989
rect 64349 118961 64383 118989
rect 64411 118961 79557 118989
rect 79585 118961 79619 118989
rect 79647 118961 79681 118989
rect 79709 118961 79743 118989
rect 79771 118961 94917 118989
rect 94945 118961 94979 118989
rect 95007 118961 95041 118989
rect 95069 118961 95103 118989
rect 95131 118961 102259 118989
rect 102287 118961 102321 118989
rect 102349 118961 117619 118989
rect 117647 118961 117681 118989
rect 117709 118961 125637 118989
rect 125665 118961 125699 118989
rect 125727 118961 125761 118989
rect 125789 118961 125823 118989
rect 125851 118961 140997 118989
rect 141025 118961 141059 118989
rect 141087 118961 141121 118989
rect 141149 118961 141183 118989
rect 141211 118961 156357 118989
rect 156385 118961 156419 118989
rect 156447 118961 156481 118989
rect 156509 118961 156543 118989
rect 156571 118961 162259 118989
rect 162287 118961 162321 118989
rect 162349 118961 177619 118989
rect 177647 118961 177681 118989
rect 177709 118961 192979 118989
rect 193007 118961 193041 118989
rect 193069 118961 208339 118989
rect 208367 118961 208401 118989
rect 208429 118961 223699 118989
rect 223727 118961 223761 118989
rect 223789 118961 239059 118989
rect 239087 118961 239121 118989
rect 239149 118961 254419 118989
rect 254447 118961 254481 118989
rect 254509 118961 269779 118989
rect 269807 118961 269841 118989
rect 269869 118961 279237 118989
rect 279265 118961 279299 118989
rect 279327 118961 279361 118989
rect 279389 118961 279423 118989
rect 279451 118961 294597 118989
rect 294625 118961 294659 118989
rect 294687 118961 294721 118989
rect 294749 118961 294783 118989
rect 294811 118961 298248 118989
rect 298276 118961 298310 118989
rect 298338 118961 298372 118989
rect 298400 118961 298434 118989
rect 298462 118961 298990 118989
rect -958 118913 298990 118961
rect -958 113175 298990 113223
rect -958 113147 -910 113175
rect -882 113147 -848 113175
rect -820 113147 -786 113175
rect -758 113147 -724 113175
rect -696 113147 4617 113175
rect 4645 113147 4679 113175
rect 4707 113147 4741 113175
rect 4769 113147 4803 113175
rect 4831 113147 19977 113175
rect 20005 113147 20039 113175
rect 20067 113147 20101 113175
rect 20129 113147 20163 113175
rect 20191 113147 35337 113175
rect 35365 113147 35399 113175
rect 35427 113147 35461 113175
rect 35489 113147 35523 113175
rect 35551 113147 50697 113175
rect 50725 113147 50759 113175
rect 50787 113147 50821 113175
rect 50849 113147 50883 113175
rect 50911 113147 66057 113175
rect 66085 113147 66119 113175
rect 66147 113147 66181 113175
rect 66209 113147 66243 113175
rect 66271 113147 81417 113175
rect 81445 113147 81479 113175
rect 81507 113147 81541 113175
rect 81569 113147 81603 113175
rect 81631 113147 96777 113175
rect 96805 113147 96839 113175
rect 96867 113147 96901 113175
rect 96929 113147 96963 113175
rect 96991 113147 109939 113175
rect 109967 113147 110001 113175
rect 110029 113147 125299 113175
rect 125327 113147 125361 113175
rect 125389 113147 127497 113175
rect 127525 113147 127559 113175
rect 127587 113147 127621 113175
rect 127649 113147 127683 113175
rect 127711 113147 142857 113175
rect 142885 113147 142919 113175
rect 142947 113147 142981 113175
rect 143009 113147 143043 113175
rect 143071 113147 158217 113175
rect 158245 113147 158279 113175
rect 158307 113147 158341 113175
rect 158369 113147 158403 113175
rect 158431 113147 169939 113175
rect 169967 113147 170001 113175
rect 170029 113147 185299 113175
rect 185327 113147 185361 113175
rect 185389 113147 200659 113175
rect 200687 113147 200721 113175
rect 200749 113147 216019 113175
rect 216047 113147 216081 113175
rect 216109 113147 231379 113175
rect 231407 113147 231441 113175
rect 231469 113147 246739 113175
rect 246767 113147 246801 113175
rect 246829 113147 262099 113175
rect 262127 113147 262161 113175
rect 262189 113147 281097 113175
rect 281125 113147 281159 113175
rect 281187 113147 281221 113175
rect 281249 113147 281283 113175
rect 281311 113147 296457 113175
rect 296485 113147 296519 113175
rect 296547 113147 296581 113175
rect 296609 113147 296643 113175
rect 296671 113147 298728 113175
rect 298756 113147 298790 113175
rect 298818 113147 298852 113175
rect 298880 113147 298914 113175
rect 298942 113147 298990 113175
rect -958 113113 298990 113147
rect -958 113085 -910 113113
rect -882 113085 -848 113113
rect -820 113085 -786 113113
rect -758 113085 -724 113113
rect -696 113085 4617 113113
rect 4645 113085 4679 113113
rect 4707 113085 4741 113113
rect 4769 113085 4803 113113
rect 4831 113085 19977 113113
rect 20005 113085 20039 113113
rect 20067 113085 20101 113113
rect 20129 113085 20163 113113
rect 20191 113085 35337 113113
rect 35365 113085 35399 113113
rect 35427 113085 35461 113113
rect 35489 113085 35523 113113
rect 35551 113085 50697 113113
rect 50725 113085 50759 113113
rect 50787 113085 50821 113113
rect 50849 113085 50883 113113
rect 50911 113085 66057 113113
rect 66085 113085 66119 113113
rect 66147 113085 66181 113113
rect 66209 113085 66243 113113
rect 66271 113085 81417 113113
rect 81445 113085 81479 113113
rect 81507 113085 81541 113113
rect 81569 113085 81603 113113
rect 81631 113085 96777 113113
rect 96805 113085 96839 113113
rect 96867 113085 96901 113113
rect 96929 113085 96963 113113
rect 96991 113085 109939 113113
rect 109967 113085 110001 113113
rect 110029 113085 125299 113113
rect 125327 113085 125361 113113
rect 125389 113085 127497 113113
rect 127525 113085 127559 113113
rect 127587 113085 127621 113113
rect 127649 113085 127683 113113
rect 127711 113085 142857 113113
rect 142885 113085 142919 113113
rect 142947 113085 142981 113113
rect 143009 113085 143043 113113
rect 143071 113085 158217 113113
rect 158245 113085 158279 113113
rect 158307 113085 158341 113113
rect 158369 113085 158403 113113
rect 158431 113085 169939 113113
rect 169967 113085 170001 113113
rect 170029 113085 185299 113113
rect 185327 113085 185361 113113
rect 185389 113085 200659 113113
rect 200687 113085 200721 113113
rect 200749 113085 216019 113113
rect 216047 113085 216081 113113
rect 216109 113085 231379 113113
rect 231407 113085 231441 113113
rect 231469 113085 246739 113113
rect 246767 113085 246801 113113
rect 246829 113085 262099 113113
rect 262127 113085 262161 113113
rect 262189 113085 281097 113113
rect 281125 113085 281159 113113
rect 281187 113085 281221 113113
rect 281249 113085 281283 113113
rect 281311 113085 296457 113113
rect 296485 113085 296519 113113
rect 296547 113085 296581 113113
rect 296609 113085 296643 113113
rect 296671 113085 298728 113113
rect 298756 113085 298790 113113
rect 298818 113085 298852 113113
rect 298880 113085 298914 113113
rect 298942 113085 298990 113113
rect -958 113051 298990 113085
rect -958 113023 -910 113051
rect -882 113023 -848 113051
rect -820 113023 -786 113051
rect -758 113023 -724 113051
rect -696 113023 4617 113051
rect 4645 113023 4679 113051
rect 4707 113023 4741 113051
rect 4769 113023 4803 113051
rect 4831 113023 19977 113051
rect 20005 113023 20039 113051
rect 20067 113023 20101 113051
rect 20129 113023 20163 113051
rect 20191 113023 35337 113051
rect 35365 113023 35399 113051
rect 35427 113023 35461 113051
rect 35489 113023 35523 113051
rect 35551 113023 50697 113051
rect 50725 113023 50759 113051
rect 50787 113023 50821 113051
rect 50849 113023 50883 113051
rect 50911 113023 66057 113051
rect 66085 113023 66119 113051
rect 66147 113023 66181 113051
rect 66209 113023 66243 113051
rect 66271 113023 81417 113051
rect 81445 113023 81479 113051
rect 81507 113023 81541 113051
rect 81569 113023 81603 113051
rect 81631 113023 96777 113051
rect 96805 113023 96839 113051
rect 96867 113023 96901 113051
rect 96929 113023 96963 113051
rect 96991 113023 109939 113051
rect 109967 113023 110001 113051
rect 110029 113023 125299 113051
rect 125327 113023 125361 113051
rect 125389 113023 127497 113051
rect 127525 113023 127559 113051
rect 127587 113023 127621 113051
rect 127649 113023 127683 113051
rect 127711 113023 142857 113051
rect 142885 113023 142919 113051
rect 142947 113023 142981 113051
rect 143009 113023 143043 113051
rect 143071 113023 158217 113051
rect 158245 113023 158279 113051
rect 158307 113023 158341 113051
rect 158369 113023 158403 113051
rect 158431 113023 169939 113051
rect 169967 113023 170001 113051
rect 170029 113023 185299 113051
rect 185327 113023 185361 113051
rect 185389 113023 200659 113051
rect 200687 113023 200721 113051
rect 200749 113023 216019 113051
rect 216047 113023 216081 113051
rect 216109 113023 231379 113051
rect 231407 113023 231441 113051
rect 231469 113023 246739 113051
rect 246767 113023 246801 113051
rect 246829 113023 262099 113051
rect 262127 113023 262161 113051
rect 262189 113023 281097 113051
rect 281125 113023 281159 113051
rect 281187 113023 281221 113051
rect 281249 113023 281283 113051
rect 281311 113023 296457 113051
rect 296485 113023 296519 113051
rect 296547 113023 296581 113051
rect 296609 113023 296643 113051
rect 296671 113023 298728 113051
rect 298756 113023 298790 113051
rect 298818 113023 298852 113051
rect 298880 113023 298914 113051
rect 298942 113023 298990 113051
rect -958 112989 298990 113023
rect -958 112961 -910 112989
rect -882 112961 -848 112989
rect -820 112961 -786 112989
rect -758 112961 -724 112989
rect -696 112961 4617 112989
rect 4645 112961 4679 112989
rect 4707 112961 4741 112989
rect 4769 112961 4803 112989
rect 4831 112961 19977 112989
rect 20005 112961 20039 112989
rect 20067 112961 20101 112989
rect 20129 112961 20163 112989
rect 20191 112961 35337 112989
rect 35365 112961 35399 112989
rect 35427 112961 35461 112989
rect 35489 112961 35523 112989
rect 35551 112961 50697 112989
rect 50725 112961 50759 112989
rect 50787 112961 50821 112989
rect 50849 112961 50883 112989
rect 50911 112961 66057 112989
rect 66085 112961 66119 112989
rect 66147 112961 66181 112989
rect 66209 112961 66243 112989
rect 66271 112961 81417 112989
rect 81445 112961 81479 112989
rect 81507 112961 81541 112989
rect 81569 112961 81603 112989
rect 81631 112961 96777 112989
rect 96805 112961 96839 112989
rect 96867 112961 96901 112989
rect 96929 112961 96963 112989
rect 96991 112961 109939 112989
rect 109967 112961 110001 112989
rect 110029 112961 125299 112989
rect 125327 112961 125361 112989
rect 125389 112961 127497 112989
rect 127525 112961 127559 112989
rect 127587 112961 127621 112989
rect 127649 112961 127683 112989
rect 127711 112961 142857 112989
rect 142885 112961 142919 112989
rect 142947 112961 142981 112989
rect 143009 112961 143043 112989
rect 143071 112961 158217 112989
rect 158245 112961 158279 112989
rect 158307 112961 158341 112989
rect 158369 112961 158403 112989
rect 158431 112961 169939 112989
rect 169967 112961 170001 112989
rect 170029 112961 185299 112989
rect 185327 112961 185361 112989
rect 185389 112961 200659 112989
rect 200687 112961 200721 112989
rect 200749 112961 216019 112989
rect 216047 112961 216081 112989
rect 216109 112961 231379 112989
rect 231407 112961 231441 112989
rect 231469 112961 246739 112989
rect 246767 112961 246801 112989
rect 246829 112961 262099 112989
rect 262127 112961 262161 112989
rect 262189 112961 281097 112989
rect 281125 112961 281159 112989
rect 281187 112961 281221 112989
rect 281249 112961 281283 112989
rect 281311 112961 296457 112989
rect 296485 112961 296519 112989
rect 296547 112961 296581 112989
rect 296609 112961 296643 112989
rect 296671 112961 298728 112989
rect 298756 112961 298790 112989
rect 298818 112961 298852 112989
rect 298880 112961 298914 112989
rect 298942 112961 298990 112989
rect -958 112913 298990 112961
rect -958 110175 298990 110223
rect -958 110147 -430 110175
rect -402 110147 -368 110175
rect -340 110147 -306 110175
rect -278 110147 -244 110175
rect -216 110147 2757 110175
rect 2785 110147 2819 110175
rect 2847 110147 2881 110175
rect 2909 110147 2943 110175
rect 2971 110147 18117 110175
rect 18145 110147 18179 110175
rect 18207 110147 18241 110175
rect 18269 110147 18303 110175
rect 18331 110147 33477 110175
rect 33505 110147 33539 110175
rect 33567 110147 33601 110175
rect 33629 110147 33663 110175
rect 33691 110147 48837 110175
rect 48865 110147 48899 110175
rect 48927 110147 48961 110175
rect 48989 110147 49023 110175
rect 49051 110147 64197 110175
rect 64225 110147 64259 110175
rect 64287 110147 64321 110175
rect 64349 110147 64383 110175
rect 64411 110147 79557 110175
rect 79585 110147 79619 110175
rect 79647 110147 79681 110175
rect 79709 110147 79743 110175
rect 79771 110147 94917 110175
rect 94945 110147 94979 110175
rect 95007 110147 95041 110175
rect 95069 110147 95103 110175
rect 95131 110147 102259 110175
rect 102287 110147 102321 110175
rect 102349 110147 117619 110175
rect 117647 110147 117681 110175
rect 117709 110147 125637 110175
rect 125665 110147 125699 110175
rect 125727 110147 125761 110175
rect 125789 110147 125823 110175
rect 125851 110147 140997 110175
rect 141025 110147 141059 110175
rect 141087 110147 141121 110175
rect 141149 110147 141183 110175
rect 141211 110147 156357 110175
rect 156385 110147 156419 110175
rect 156447 110147 156481 110175
rect 156509 110147 156543 110175
rect 156571 110147 162259 110175
rect 162287 110147 162321 110175
rect 162349 110147 177619 110175
rect 177647 110147 177681 110175
rect 177709 110147 192979 110175
rect 193007 110147 193041 110175
rect 193069 110147 208339 110175
rect 208367 110147 208401 110175
rect 208429 110147 223699 110175
rect 223727 110147 223761 110175
rect 223789 110147 239059 110175
rect 239087 110147 239121 110175
rect 239149 110147 254419 110175
rect 254447 110147 254481 110175
rect 254509 110147 269779 110175
rect 269807 110147 269841 110175
rect 269869 110147 279237 110175
rect 279265 110147 279299 110175
rect 279327 110147 279361 110175
rect 279389 110147 279423 110175
rect 279451 110147 294597 110175
rect 294625 110147 294659 110175
rect 294687 110147 294721 110175
rect 294749 110147 294783 110175
rect 294811 110147 298248 110175
rect 298276 110147 298310 110175
rect 298338 110147 298372 110175
rect 298400 110147 298434 110175
rect 298462 110147 298990 110175
rect -958 110113 298990 110147
rect -958 110085 -430 110113
rect -402 110085 -368 110113
rect -340 110085 -306 110113
rect -278 110085 -244 110113
rect -216 110085 2757 110113
rect 2785 110085 2819 110113
rect 2847 110085 2881 110113
rect 2909 110085 2943 110113
rect 2971 110085 18117 110113
rect 18145 110085 18179 110113
rect 18207 110085 18241 110113
rect 18269 110085 18303 110113
rect 18331 110085 33477 110113
rect 33505 110085 33539 110113
rect 33567 110085 33601 110113
rect 33629 110085 33663 110113
rect 33691 110085 48837 110113
rect 48865 110085 48899 110113
rect 48927 110085 48961 110113
rect 48989 110085 49023 110113
rect 49051 110085 64197 110113
rect 64225 110085 64259 110113
rect 64287 110085 64321 110113
rect 64349 110085 64383 110113
rect 64411 110085 79557 110113
rect 79585 110085 79619 110113
rect 79647 110085 79681 110113
rect 79709 110085 79743 110113
rect 79771 110085 94917 110113
rect 94945 110085 94979 110113
rect 95007 110085 95041 110113
rect 95069 110085 95103 110113
rect 95131 110085 102259 110113
rect 102287 110085 102321 110113
rect 102349 110085 117619 110113
rect 117647 110085 117681 110113
rect 117709 110085 125637 110113
rect 125665 110085 125699 110113
rect 125727 110085 125761 110113
rect 125789 110085 125823 110113
rect 125851 110085 140997 110113
rect 141025 110085 141059 110113
rect 141087 110085 141121 110113
rect 141149 110085 141183 110113
rect 141211 110085 156357 110113
rect 156385 110085 156419 110113
rect 156447 110085 156481 110113
rect 156509 110085 156543 110113
rect 156571 110085 162259 110113
rect 162287 110085 162321 110113
rect 162349 110085 177619 110113
rect 177647 110085 177681 110113
rect 177709 110085 192979 110113
rect 193007 110085 193041 110113
rect 193069 110085 208339 110113
rect 208367 110085 208401 110113
rect 208429 110085 223699 110113
rect 223727 110085 223761 110113
rect 223789 110085 239059 110113
rect 239087 110085 239121 110113
rect 239149 110085 254419 110113
rect 254447 110085 254481 110113
rect 254509 110085 269779 110113
rect 269807 110085 269841 110113
rect 269869 110085 279237 110113
rect 279265 110085 279299 110113
rect 279327 110085 279361 110113
rect 279389 110085 279423 110113
rect 279451 110085 294597 110113
rect 294625 110085 294659 110113
rect 294687 110085 294721 110113
rect 294749 110085 294783 110113
rect 294811 110085 298248 110113
rect 298276 110085 298310 110113
rect 298338 110085 298372 110113
rect 298400 110085 298434 110113
rect 298462 110085 298990 110113
rect -958 110051 298990 110085
rect -958 110023 -430 110051
rect -402 110023 -368 110051
rect -340 110023 -306 110051
rect -278 110023 -244 110051
rect -216 110023 2757 110051
rect 2785 110023 2819 110051
rect 2847 110023 2881 110051
rect 2909 110023 2943 110051
rect 2971 110023 18117 110051
rect 18145 110023 18179 110051
rect 18207 110023 18241 110051
rect 18269 110023 18303 110051
rect 18331 110023 33477 110051
rect 33505 110023 33539 110051
rect 33567 110023 33601 110051
rect 33629 110023 33663 110051
rect 33691 110023 48837 110051
rect 48865 110023 48899 110051
rect 48927 110023 48961 110051
rect 48989 110023 49023 110051
rect 49051 110023 64197 110051
rect 64225 110023 64259 110051
rect 64287 110023 64321 110051
rect 64349 110023 64383 110051
rect 64411 110023 79557 110051
rect 79585 110023 79619 110051
rect 79647 110023 79681 110051
rect 79709 110023 79743 110051
rect 79771 110023 94917 110051
rect 94945 110023 94979 110051
rect 95007 110023 95041 110051
rect 95069 110023 95103 110051
rect 95131 110023 102259 110051
rect 102287 110023 102321 110051
rect 102349 110023 117619 110051
rect 117647 110023 117681 110051
rect 117709 110023 125637 110051
rect 125665 110023 125699 110051
rect 125727 110023 125761 110051
rect 125789 110023 125823 110051
rect 125851 110023 140997 110051
rect 141025 110023 141059 110051
rect 141087 110023 141121 110051
rect 141149 110023 141183 110051
rect 141211 110023 156357 110051
rect 156385 110023 156419 110051
rect 156447 110023 156481 110051
rect 156509 110023 156543 110051
rect 156571 110023 162259 110051
rect 162287 110023 162321 110051
rect 162349 110023 177619 110051
rect 177647 110023 177681 110051
rect 177709 110023 192979 110051
rect 193007 110023 193041 110051
rect 193069 110023 208339 110051
rect 208367 110023 208401 110051
rect 208429 110023 223699 110051
rect 223727 110023 223761 110051
rect 223789 110023 239059 110051
rect 239087 110023 239121 110051
rect 239149 110023 254419 110051
rect 254447 110023 254481 110051
rect 254509 110023 269779 110051
rect 269807 110023 269841 110051
rect 269869 110023 279237 110051
rect 279265 110023 279299 110051
rect 279327 110023 279361 110051
rect 279389 110023 279423 110051
rect 279451 110023 294597 110051
rect 294625 110023 294659 110051
rect 294687 110023 294721 110051
rect 294749 110023 294783 110051
rect 294811 110023 298248 110051
rect 298276 110023 298310 110051
rect 298338 110023 298372 110051
rect 298400 110023 298434 110051
rect 298462 110023 298990 110051
rect -958 109989 298990 110023
rect -958 109961 -430 109989
rect -402 109961 -368 109989
rect -340 109961 -306 109989
rect -278 109961 -244 109989
rect -216 109961 2757 109989
rect 2785 109961 2819 109989
rect 2847 109961 2881 109989
rect 2909 109961 2943 109989
rect 2971 109961 18117 109989
rect 18145 109961 18179 109989
rect 18207 109961 18241 109989
rect 18269 109961 18303 109989
rect 18331 109961 33477 109989
rect 33505 109961 33539 109989
rect 33567 109961 33601 109989
rect 33629 109961 33663 109989
rect 33691 109961 48837 109989
rect 48865 109961 48899 109989
rect 48927 109961 48961 109989
rect 48989 109961 49023 109989
rect 49051 109961 64197 109989
rect 64225 109961 64259 109989
rect 64287 109961 64321 109989
rect 64349 109961 64383 109989
rect 64411 109961 79557 109989
rect 79585 109961 79619 109989
rect 79647 109961 79681 109989
rect 79709 109961 79743 109989
rect 79771 109961 94917 109989
rect 94945 109961 94979 109989
rect 95007 109961 95041 109989
rect 95069 109961 95103 109989
rect 95131 109961 102259 109989
rect 102287 109961 102321 109989
rect 102349 109961 117619 109989
rect 117647 109961 117681 109989
rect 117709 109961 125637 109989
rect 125665 109961 125699 109989
rect 125727 109961 125761 109989
rect 125789 109961 125823 109989
rect 125851 109961 140997 109989
rect 141025 109961 141059 109989
rect 141087 109961 141121 109989
rect 141149 109961 141183 109989
rect 141211 109961 156357 109989
rect 156385 109961 156419 109989
rect 156447 109961 156481 109989
rect 156509 109961 156543 109989
rect 156571 109961 162259 109989
rect 162287 109961 162321 109989
rect 162349 109961 177619 109989
rect 177647 109961 177681 109989
rect 177709 109961 192979 109989
rect 193007 109961 193041 109989
rect 193069 109961 208339 109989
rect 208367 109961 208401 109989
rect 208429 109961 223699 109989
rect 223727 109961 223761 109989
rect 223789 109961 239059 109989
rect 239087 109961 239121 109989
rect 239149 109961 254419 109989
rect 254447 109961 254481 109989
rect 254509 109961 269779 109989
rect 269807 109961 269841 109989
rect 269869 109961 279237 109989
rect 279265 109961 279299 109989
rect 279327 109961 279361 109989
rect 279389 109961 279423 109989
rect 279451 109961 294597 109989
rect 294625 109961 294659 109989
rect 294687 109961 294721 109989
rect 294749 109961 294783 109989
rect 294811 109961 298248 109989
rect 298276 109961 298310 109989
rect 298338 109961 298372 109989
rect 298400 109961 298434 109989
rect 298462 109961 298990 109989
rect -958 109913 298990 109961
rect -958 104175 298990 104223
rect -958 104147 -910 104175
rect -882 104147 -848 104175
rect -820 104147 -786 104175
rect -758 104147 -724 104175
rect -696 104147 4617 104175
rect 4645 104147 4679 104175
rect 4707 104147 4741 104175
rect 4769 104147 4803 104175
rect 4831 104147 19977 104175
rect 20005 104147 20039 104175
rect 20067 104147 20101 104175
rect 20129 104147 20163 104175
rect 20191 104147 35337 104175
rect 35365 104147 35399 104175
rect 35427 104147 35461 104175
rect 35489 104147 35523 104175
rect 35551 104147 50697 104175
rect 50725 104147 50759 104175
rect 50787 104147 50821 104175
rect 50849 104147 50883 104175
rect 50911 104147 66057 104175
rect 66085 104147 66119 104175
rect 66147 104147 66181 104175
rect 66209 104147 66243 104175
rect 66271 104147 81417 104175
rect 81445 104147 81479 104175
rect 81507 104147 81541 104175
rect 81569 104147 81603 104175
rect 81631 104147 96777 104175
rect 96805 104147 96839 104175
rect 96867 104147 96901 104175
rect 96929 104147 96963 104175
rect 96991 104147 109939 104175
rect 109967 104147 110001 104175
rect 110029 104147 125299 104175
rect 125327 104147 125361 104175
rect 125389 104147 127497 104175
rect 127525 104147 127559 104175
rect 127587 104147 127621 104175
rect 127649 104147 127683 104175
rect 127711 104147 142857 104175
rect 142885 104147 142919 104175
rect 142947 104147 142981 104175
rect 143009 104147 143043 104175
rect 143071 104147 158217 104175
rect 158245 104147 158279 104175
rect 158307 104147 158341 104175
rect 158369 104147 158403 104175
rect 158431 104147 169939 104175
rect 169967 104147 170001 104175
rect 170029 104147 185299 104175
rect 185327 104147 185361 104175
rect 185389 104147 200659 104175
rect 200687 104147 200721 104175
rect 200749 104147 216019 104175
rect 216047 104147 216081 104175
rect 216109 104147 231379 104175
rect 231407 104147 231441 104175
rect 231469 104147 246739 104175
rect 246767 104147 246801 104175
rect 246829 104147 262099 104175
rect 262127 104147 262161 104175
rect 262189 104147 281097 104175
rect 281125 104147 281159 104175
rect 281187 104147 281221 104175
rect 281249 104147 281283 104175
rect 281311 104147 296457 104175
rect 296485 104147 296519 104175
rect 296547 104147 296581 104175
rect 296609 104147 296643 104175
rect 296671 104147 298728 104175
rect 298756 104147 298790 104175
rect 298818 104147 298852 104175
rect 298880 104147 298914 104175
rect 298942 104147 298990 104175
rect -958 104113 298990 104147
rect -958 104085 -910 104113
rect -882 104085 -848 104113
rect -820 104085 -786 104113
rect -758 104085 -724 104113
rect -696 104085 4617 104113
rect 4645 104085 4679 104113
rect 4707 104085 4741 104113
rect 4769 104085 4803 104113
rect 4831 104085 19977 104113
rect 20005 104085 20039 104113
rect 20067 104085 20101 104113
rect 20129 104085 20163 104113
rect 20191 104085 35337 104113
rect 35365 104085 35399 104113
rect 35427 104085 35461 104113
rect 35489 104085 35523 104113
rect 35551 104085 50697 104113
rect 50725 104085 50759 104113
rect 50787 104085 50821 104113
rect 50849 104085 50883 104113
rect 50911 104085 66057 104113
rect 66085 104085 66119 104113
rect 66147 104085 66181 104113
rect 66209 104085 66243 104113
rect 66271 104085 81417 104113
rect 81445 104085 81479 104113
rect 81507 104085 81541 104113
rect 81569 104085 81603 104113
rect 81631 104085 96777 104113
rect 96805 104085 96839 104113
rect 96867 104085 96901 104113
rect 96929 104085 96963 104113
rect 96991 104085 109939 104113
rect 109967 104085 110001 104113
rect 110029 104085 125299 104113
rect 125327 104085 125361 104113
rect 125389 104085 127497 104113
rect 127525 104085 127559 104113
rect 127587 104085 127621 104113
rect 127649 104085 127683 104113
rect 127711 104085 142857 104113
rect 142885 104085 142919 104113
rect 142947 104085 142981 104113
rect 143009 104085 143043 104113
rect 143071 104085 158217 104113
rect 158245 104085 158279 104113
rect 158307 104085 158341 104113
rect 158369 104085 158403 104113
rect 158431 104085 169939 104113
rect 169967 104085 170001 104113
rect 170029 104085 185299 104113
rect 185327 104085 185361 104113
rect 185389 104085 200659 104113
rect 200687 104085 200721 104113
rect 200749 104085 216019 104113
rect 216047 104085 216081 104113
rect 216109 104085 231379 104113
rect 231407 104085 231441 104113
rect 231469 104085 246739 104113
rect 246767 104085 246801 104113
rect 246829 104085 262099 104113
rect 262127 104085 262161 104113
rect 262189 104085 281097 104113
rect 281125 104085 281159 104113
rect 281187 104085 281221 104113
rect 281249 104085 281283 104113
rect 281311 104085 296457 104113
rect 296485 104085 296519 104113
rect 296547 104085 296581 104113
rect 296609 104085 296643 104113
rect 296671 104085 298728 104113
rect 298756 104085 298790 104113
rect 298818 104085 298852 104113
rect 298880 104085 298914 104113
rect 298942 104085 298990 104113
rect -958 104051 298990 104085
rect -958 104023 -910 104051
rect -882 104023 -848 104051
rect -820 104023 -786 104051
rect -758 104023 -724 104051
rect -696 104023 4617 104051
rect 4645 104023 4679 104051
rect 4707 104023 4741 104051
rect 4769 104023 4803 104051
rect 4831 104023 19977 104051
rect 20005 104023 20039 104051
rect 20067 104023 20101 104051
rect 20129 104023 20163 104051
rect 20191 104023 35337 104051
rect 35365 104023 35399 104051
rect 35427 104023 35461 104051
rect 35489 104023 35523 104051
rect 35551 104023 50697 104051
rect 50725 104023 50759 104051
rect 50787 104023 50821 104051
rect 50849 104023 50883 104051
rect 50911 104023 66057 104051
rect 66085 104023 66119 104051
rect 66147 104023 66181 104051
rect 66209 104023 66243 104051
rect 66271 104023 81417 104051
rect 81445 104023 81479 104051
rect 81507 104023 81541 104051
rect 81569 104023 81603 104051
rect 81631 104023 96777 104051
rect 96805 104023 96839 104051
rect 96867 104023 96901 104051
rect 96929 104023 96963 104051
rect 96991 104023 109939 104051
rect 109967 104023 110001 104051
rect 110029 104023 125299 104051
rect 125327 104023 125361 104051
rect 125389 104023 127497 104051
rect 127525 104023 127559 104051
rect 127587 104023 127621 104051
rect 127649 104023 127683 104051
rect 127711 104023 142857 104051
rect 142885 104023 142919 104051
rect 142947 104023 142981 104051
rect 143009 104023 143043 104051
rect 143071 104023 158217 104051
rect 158245 104023 158279 104051
rect 158307 104023 158341 104051
rect 158369 104023 158403 104051
rect 158431 104023 169939 104051
rect 169967 104023 170001 104051
rect 170029 104023 185299 104051
rect 185327 104023 185361 104051
rect 185389 104023 200659 104051
rect 200687 104023 200721 104051
rect 200749 104023 216019 104051
rect 216047 104023 216081 104051
rect 216109 104023 231379 104051
rect 231407 104023 231441 104051
rect 231469 104023 246739 104051
rect 246767 104023 246801 104051
rect 246829 104023 262099 104051
rect 262127 104023 262161 104051
rect 262189 104023 281097 104051
rect 281125 104023 281159 104051
rect 281187 104023 281221 104051
rect 281249 104023 281283 104051
rect 281311 104023 296457 104051
rect 296485 104023 296519 104051
rect 296547 104023 296581 104051
rect 296609 104023 296643 104051
rect 296671 104023 298728 104051
rect 298756 104023 298790 104051
rect 298818 104023 298852 104051
rect 298880 104023 298914 104051
rect 298942 104023 298990 104051
rect -958 103989 298990 104023
rect -958 103961 -910 103989
rect -882 103961 -848 103989
rect -820 103961 -786 103989
rect -758 103961 -724 103989
rect -696 103961 4617 103989
rect 4645 103961 4679 103989
rect 4707 103961 4741 103989
rect 4769 103961 4803 103989
rect 4831 103961 19977 103989
rect 20005 103961 20039 103989
rect 20067 103961 20101 103989
rect 20129 103961 20163 103989
rect 20191 103961 35337 103989
rect 35365 103961 35399 103989
rect 35427 103961 35461 103989
rect 35489 103961 35523 103989
rect 35551 103961 50697 103989
rect 50725 103961 50759 103989
rect 50787 103961 50821 103989
rect 50849 103961 50883 103989
rect 50911 103961 66057 103989
rect 66085 103961 66119 103989
rect 66147 103961 66181 103989
rect 66209 103961 66243 103989
rect 66271 103961 81417 103989
rect 81445 103961 81479 103989
rect 81507 103961 81541 103989
rect 81569 103961 81603 103989
rect 81631 103961 96777 103989
rect 96805 103961 96839 103989
rect 96867 103961 96901 103989
rect 96929 103961 96963 103989
rect 96991 103961 109939 103989
rect 109967 103961 110001 103989
rect 110029 103961 125299 103989
rect 125327 103961 125361 103989
rect 125389 103961 127497 103989
rect 127525 103961 127559 103989
rect 127587 103961 127621 103989
rect 127649 103961 127683 103989
rect 127711 103961 142857 103989
rect 142885 103961 142919 103989
rect 142947 103961 142981 103989
rect 143009 103961 143043 103989
rect 143071 103961 158217 103989
rect 158245 103961 158279 103989
rect 158307 103961 158341 103989
rect 158369 103961 158403 103989
rect 158431 103961 169939 103989
rect 169967 103961 170001 103989
rect 170029 103961 185299 103989
rect 185327 103961 185361 103989
rect 185389 103961 200659 103989
rect 200687 103961 200721 103989
rect 200749 103961 216019 103989
rect 216047 103961 216081 103989
rect 216109 103961 231379 103989
rect 231407 103961 231441 103989
rect 231469 103961 246739 103989
rect 246767 103961 246801 103989
rect 246829 103961 262099 103989
rect 262127 103961 262161 103989
rect 262189 103961 281097 103989
rect 281125 103961 281159 103989
rect 281187 103961 281221 103989
rect 281249 103961 281283 103989
rect 281311 103961 296457 103989
rect 296485 103961 296519 103989
rect 296547 103961 296581 103989
rect 296609 103961 296643 103989
rect 296671 103961 298728 103989
rect 298756 103961 298790 103989
rect 298818 103961 298852 103989
rect 298880 103961 298914 103989
rect 298942 103961 298990 103989
rect -958 103913 298990 103961
rect -958 101175 298990 101223
rect -958 101147 -430 101175
rect -402 101147 -368 101175
rect -340 101147 -306 101175
rect -278 101147 -244 101175
rect -216 101147 2757 101175
rect 2785 101147 2819 101175
rect 2847 101147 2881 101175
rect 2909 101147 2943 101175
rect 2971 101147 16259 101175
rect 16287 101147 16321 101175
rect 16349 101147 18117 101175
rect 18145 101147 18179 101175
rect 18207 101147 18241 101175
rect 18269 101147 18303 101175
rect 18331 101147 31619 101175
rect 31647 101147 31681 101175
rect 31709 101147 33477 101175
rect 33505 101147 33539 101175
rect 33567 101147 33601 101175
rect 33629 101147 33663 101175
rect 33691 101147 46979 101175
rect 47007 101147 47041 101175
rect 47069 101147 48837 101175
rect 48865 101147 48899 101175
rect 48927 101147 48961 101175
rect 48989 101147 49023 101175
rect 49051 101147 62339 101175
rect 62367 101147 62401 101175
rect 62429 101147 64197 101175
rect 64225 101147 64259 101175
rect 64287 101147 64321 101175
rect 64349 101147 64383 101175
rect 64411 101147 77699 101175
rect 77727 101147 77761 101175
rect 77789 101147 79557 101175
rect 79585 101147 79619 101175
rect 79647 101147 79681 101175
rect 79709 101147 79743 101175
rect 79771 101147 93059 101175
rect 93087 101147 93121 101175
rect 93149 101147 94917 101175
rect 94945 101147 94979 101175
rect 95007 101147 95041 101175
rect 95069 101147 95103 101175
rect 95131 101147 102259 101175
rect 102287 101147 102321 101175
rect 102349 101147 117619 101175
rect 117647 101147 117681 101175
rect 117709 101147 125637 101175
rect 125665 101147 125699 101175
rect 125727 101147 125761 101175
rect 125789 101147 125823 101175
rect 125851 101147 140997 101175
rect 141025 101147 141059 101175
rect 141087 101147 141121 101175
rect 141149 101147 141183 101175
rect 141211 101147 156357 101175
rect 156385 101147 156419 101175
rect 156447 101147 156481 101175
rect 156509 101147 156543 101175
rect 156571 101147 162259 101175
rect 162287 101147 162321 101175
rect 162349 101147 177619 101175
rect 177647 101147 177681 101175
rect 177709 101147 192979 101175
rect 193007 101147 193041 101175
rect 193069 101147 208339 101175
rect 208367 101147 208401 101175
rect 208429 101147 223699 101175
rect 223727 101147 223761 101175
rect 223789 101147 239059 101175
rect 239087 101147 239121 101175
rect 239149 101147 254419 101175
rect 254447 101147 254481 101175
rect 254509 101147 269779 101175
rect 269807 101147 269841 101175
rect 269869 101147 279237 101175
rect 279265 101147 279299 101175
rect 279327 101147 279361 101175
rect 279389 101147 279423 101175
rect 279451 101147 294597 101175
rect 294625 101147 294659 101175
rect 294687 101147 294721 101175
rect 294749 101147 294783 101175
rect 294811 101147 298248 101175
rect 298276 101147 298310 101175
rect 298338 101147 298372 101175
rect 298400 101147 298434 101175
rect 298462 101147 298990 101175
rect -958 101113 298990 101147
rect -958 101085 -430 101113
rect -402 101085 -368 101113
rect -340 101085 -306 101113
rect -278 101085 -244 101113
rect -216 101085 2757 101113
rect 2785 101085 2819 101113
rect 2847 101085 2881 101113
rect 2909 101085 2943 101113
rect 2971 101085 16259 101113
rect 16287 101085 16321 101113
rect 16349 101085 18117 101113
rect 18145 101085 18179 101113
rect 18207 101085 18241 101113
rect 18269 101085 18303 101113
rect 18331 101085 31619 101113
rect 31647 101085 31681 101113
rect 31709 101085 33477 101113
rect 33505 101085 33539 101113
rect 33567 101085 33601 101113
rect 33629 101085 33663 101113
rect 33691 101085 46979 101113
rect 47007 101085 47041 101113
rect 47069 101085 48837 101113
rect 48865 101085 48899 101113
rect 48927 101085 48961 101113
rect 48989 101085 49023 101113
rect 49051 101085 62339 101113
rect 62367 101085 62401 101113
rect 62429 101085 64197 101113
rect 64225 101085 64259 101113
rect 64287 101085 64321 101113
rect 64349 101085 64383 101113
rect 64411 101085 77699 101113
rect 77727 101085 77761 101113
rect 77789 101085 79557 101113
rect 79585 101085 79619 101113
rect 79647 101085 79681 101113
rect 79709 101085 79743 101113
rect 79771 101085 93059 101113
rect 93087 101085 93121 101113
rect 93149 101085 94917 101113
rect 94945 101085 94979 101113
rect 95007 101085 95041 101113
rect 95069 101085 95103 101113
rect 95131 101085 102259 101113
rect 102287 101085 102321 101113
rect 102349 101085 117619 101113
rect 117647 101085 117681 101113
rect 117709 101085 125637 101113
rect 125665 101085 125699 101113
rect 125727 101085 125761 101113
rect 125789 101085 125823 101113
rect 125851 101085 140997 101113
rect 141025 101085 141059 101113
rect 141087 101085 141121 101113
rect 141149 101085 141183 101113
rect 141211 101085 156357 101113
rect 156385 101085 156419 101113
rect 156447 101085 156481 101113
rect 156509 101085 156543 101113
rect 156571 101085 162259 101113
rect 162287 101085 162321 101113
rect 162349 101085 177619 101113
rect 177647 101085 177681 101113
rect 177709 101085 192979 101113
rect 193007 101085 193041 101113
rect 193069 101085 208339 101113
rect 208367 101085 208401 101113
rect 208429 101085 223699 101113
rect 223727 101085 223761 101113
rect 223789 101085 239059 101113
rect 239087 101085 239121 101113
rect 239149 101085 254419 101113
rect 254447 101085 254481 101113
rect 254509 101085 269779 101113
rect 269807 101085 269841 101113
rect 269869 101085 279237 101113
rect 279265 101085 279299 101113
rect 279327 101085 279361 101113
rect 279389 101085 279423 101113
rect 279451 101085 294597 101113
rect 294625 101085 294659 101113
rect 294687 101085 294721 101113
rect 294749 101085 294783 101113
rect 294811 101085 298248 101113
rect 298276 101085 298310 101113
rect 298338 101085 298372 101113
rect 298400 101085 298434 101113
rect 298462 101085 298990 101113
rect -958 101051 298990 101085
rect -958 101023 -430 101051
rect -402 101023 -368 101051
rect -340 101023 -306 101051
rect -278 101023 -244 101051
rect -216 101023 2757 101051
rect 2785 101023 2819 101051
rect 2847 101023 2881 101051
rect 2909 101023 2943 101051
rect 2971 101023 16259 101051
rect 16287 101023 16321 101051
rect 16349 101023 18117 101051
rect 18145 101023 18179 101051
rect 18207 101023 18241 101051
rect 18269 101023 18303 101051
rect 18331 101023 31619 101051
rect 31647 101023 31681 101051
rect 31709 101023 33477 101051
rect 33505 101023 33539 101051
rect 33567 101023 33601 101051
rect 33629 101023 33663 101051
rect 33691 101023 46979 101051
rect 47007 101023 47041 101051
rect 47069 101023 48837 101051
rect 48865 101023 48899 101051
rect 48927 101023 48961 101051
rect 48989 101023 49023 101051
rect 49051 101023 62339 101051
rect 62367 101023 62401 101051
rect 62429 101023 64197 101051
rect 64225 101023 64259 101051
rect 64287 101023 64321 101051
rect 64349 101023 64383 101051
rect 64411 101023 77699 101051
rect 77727 101023 77761 101051
rect 77789 101023 79557 101051
rect 79585 101023 79619 101051
rect 79647 101023 79681 101051
rect 79709 101023 79743 101051
rect 79771 101023 93059 101051
rect 93087 101023 93121 101051
rect 93149 101023 94917 101051
rect 94945 101023 94979 101051
rect 95007 101023 95041 101051
rect 95069 101023 95103 101051
rect 95131 101023 102259 101051
rect 102287 101023 102321 101051
rect 102349 101023 117619 101051
rect 117647 101023 117681 101051
rect 117709 101023 125637 101051
rect 125665 101023 125699 101051
rect 125727 101023 125761 101051
rect 125789 101023 125823 101051
rect 125851 101023 140997 101051
rect 141025 101023 141059 101051
rect 141087 101023 141121 101051
rect 141149 101023 141183 101051
rect 141211 101023 156357 101051
rect 156385 101023 156419 101051
rect 156447 101023 156481 101051
rect 156509 101023 156543 101051
rect 156571 101023 162259 101051
rect 162287 101023 162321 101051
rect 162349 101023 177619 101051
rect 177647 101023 177681 101051
rect 177709 101023 192979 101051
rect 193007 101023 193041 101051
rect 193069 101023 208339 101051
rect 208367 101023 208401 101051
rect 208429 101023 223699 101051
rect 223727 101023 223761 101051
rect 223789 101023 239059 101051
rect 239087 101023 239121 101051
rect 239149 101023 254419 101051
rect 254447 101023 254481 101051
rect 254509 101023 269779 101051
rect 269807 101023 269841 101051
rect 269869 101023 279237 101051
rect 279265 101023 279299 101051
rect 279327 101023 279361 101051
rect 279389 101023 279423 101051
rect 279451 101023 294597 101051
rect 294625 101023 294659 101051
rect 294687 101023 294721 101051
rect 294749 101023 294783 101051
rect 294811 101023 298248 101051
rect 298276 101023 298310 101051
rect 298338 101023 298372 101051
rect 298400 101023 298434 101051
rect 298462 101023 298990 101051
rect -958 100989 298990 101023
rect -958 100961 -430 100989
rect -402 100961 -368 100989
rect -340 100961 -306 100989
rect -278 100961 -244 100989
rect -216 100961 2757 100989
rect 2785 100961 2819 100989
rect 2847 100961 2881 100989
rect 2909 100961 2943 100989
rect 2971 100961 16259 100989
rect 16287 100961 16321 100989
rect 16349 100961 18117 100989
rect 18145 100961 18179 100989
rect 18207 100961 18241 100989
rect 18269 100961 18303 100989
rect 18331 100961 31619 100989
rect 31647 100961 31681 100989
rect 31709 100961 33477 100989
rect 33505 100961 33539 100989
rect 33567 100961 33601 100989
rect 33629 100961 33663 100989
rect 33691 100961 46979 100989
rect 47007 100961 47041 100989
rect 47069 100961 48837 100989
rect 48865 100961 48899 100989
rect 48927 100961 48961 100989
rect 48989 100961 49023 100989
rect 49051 100961 62339 100989
rect 62367 100961 62401 100989
rect 62429 100961 64197 100989
rect 64225 100961 64259 100989
rect 64287 100961 64321 100989
rect 64349 100961 64383 100989
rect 64411 100961 77699 100989
rect 77727 100961 77761 100989
rect 77789 100961 79557 100989
rect 79585 100961 79619 100989
rect 79647 100961 79681 100989
rect 79709 100961 79743 100989
rect 79771 100961 93059 100989
rect 93087 100961 93121 100989
rect 93149 100961 94917 100989
rect 94945 100961 94979 100989
rect 95007 100961 95041 100989
rect 95069 100961 95103 100989
rect 95131 100961 102259 100989
rect 102287 100961 102321 100989
rect 102349 100961 117619 100989
rect 117647 100961 117681 100989
rect 117709 100961 125637 100989
rect 125665 100961 125699 100989
rect 125727 100961 125761 100989
rect 125789 100961 125823 100989
rect 125851 100961 140997 100989
rect 141025 100961 141059 100989
rect 141087 100961 141121 100989
rect 141149 100961 141183 100989
rect 141211 100961 156357 100989
rect 156385 100961 156419 100989
rect 156447 100961 156481 100989
rect 156509 100961 156543 100989
rect 156571 100961 162259 100989
rect 162287 100961 162321 100989
rect 162349 100961 177619 100989
rect 177647 100961 177681 100989
rect 177709 100961 192979 100989
rect 193007 100961 193041 100989
rect 193069 100961 208339 100989
rect 208367 100961 208401 100989
rect 208429 100961 223699 100989
rect 223727 100961 223761 100989
rect 223789 100961 239059 100989
rect 239087 100961 239121 100989
rect 239149 100961 254419 100989
rect 254447 100961 254481 100989
rect 254509 100961 269779 100989
rect 269807 100961 269841 100989
rect 269869 100961 279237 100989
rect 279265 100961 279299 100989
rect 279327 100961 279361 100989
rect 279389 100961 279423 100989
rect 279451 100961 294597 100989
rect 294625 100961 294659 100989
rect 294687 100961 294721 100989
rect 294749 100961 294783 100989
rect 294811 100961 298248 100989
rect 298276 100961 298310 100989
rect 298338 100961 298372 100989
rect 298400 100961 298434 100989
rect 298462 100961 298990 100989
rect -958 100913 298990 100961
rect -958 95175 298990 95223
rect -958 95147 -910 95175
rect -882 95147 -848 95175
rect -820 95147 -786 95175
rect -758 95147 -724 95175
rect -696 95147 4617 95175
rect 4645 95147 4679 95175
rect 4707 95147 4741 95175
rect 4769 95147 4803 95175
rect 4831 95147 19977 95175
rect 20005 95147 20039 95175
rect 20067 95147 20101 95175
rect 20129 95147 20163 95175
rect 20191 95147 23939 95175
rect 23967 95147 24001 95175
rect 24029 95147 35337 95175
rect 35365 95147 35399 95175
rect 35427 95147 35461 95175
rect 35489 95147 35523 95175
rect 35551 95147 39299 95175
rect 39327 95147 39361 95175
rect 39389 95147 50697 95175
rect 50725 95147 50759 95175
rect 50787 95147 50821 95175
rect 50849 95147 50883 95175
rect 50911 95147 54659 95175
rect 54687 95147 54721 95175
rect 54749 95147 66057 95175
rect 66085 95147 66119 95175
rect 66147 95147 66181 95175
rect 66209 95147 66243 95175
rect 66271 95147 70019 95175
rect 70047 95147 70081 95175
rect 70109 95147 81417 95175
rect 81445 95147 81479 95175
rect 81507 95147 81541 95175
rect 81569 95147 81603 95175
rect 81631 95147 85379 95175
rect 85407 95147 85441 95175
rect 85469 95147 96777 95175
rect 96805 95147 96839 95175
rect 96867 95147 96901 95175
rect 96929 95147 96963 95175
rect 96991 95147 112137 95175
rect 112165 95147 112199 95175
rect 112227 95147 112261 95175
rect 112289 95147 112323 95175
rect 112351 95147 127497 95175
rect 127525 95147 127559 95175
rect 127587 95147 127621 95175
rect 127649 95147 127683 95175
rect 127711 95147 142857 95175
rect 142885 95147 142919 95175
rect 142947 95147 142981 95175
rect 143009 95147 143043 95175
rect 143071 95147 158217 95175
rect 158245 95147 158279 95175
rect 158307 95147 158341 95175
rect 158369 95147 158403 95175
rect 158431 95147 169939 95175
rect 169967 95147 170001 95175
rect 170029 95147 185299 95175
rect 185327 95147 185361 95175
rect 185389 95147 200659 95175
rect 200687 95147 200721 95175
rect 200749 95147 216019 95175
rect 216047 95147 216081 95175
rect 216109 95147 231379 95175
rect 231407 95147 231441 95175
rect 231469 95147 246739 95175
rect 246767 95147 246801 95175
rect 246829 95147 262099 95175
rect 262127 95147 262161 95175
rect 262189 95147 281097 95175
rect 281125 95147 281159 95175
rect 281187 95147 281221 95175
rect 281249 95147 281283 95175
rect 281311 95147 296457 95175
rect 296485 95147 296519 95175
rect 296547 95147 296581 95175
rect 296609 95147 296643 95175
rect 296671 95147 298728 95175
rect 298756 95147 298790 95175
rect 298818 95147 298852 95175
rect 298880 95147 298914 95175
rect 298942 95147 298990 95175
rect -958 95113 298990 95147
rect -958 95085 -910 95113
rect -882 95085 -848 95113
rect -820 95085 -786 95113
rect -758 95085 -724 95113
rect -696 95085 4617 95113
rect 4645 95085 4679 95113
rect 4707 95085 4741 95113
rect 4769 95085 4803 95113
rect 4831 95085 19977 95113
rect 20005 95085 20039 95113
rect 20067 95085 20101 95113
rect 20129 95085 20163 95113
rect 20191 95085 23939 95113
rect 23967 95085 24001 95113
rect 24029 95085 35337 95113
rect 35365 95085 35399 95113
rect 35427 95085 35461 95113
rect 35489 95085 35523 95113
rect 35551 95085 39299 95113
rect 39327 95085 39361 95113
rect 39389 95085 50697 95113
rect 50725 95085 50759 95113
rect 50787 95085 50821 95113
rect 50849 95085 50883 95113
rect 50911 95085 54659 95113
rect 54687 95085 54721 95113
rect 54749 95085 66057 95113
rect 66085 95085 66119 95113
rect 66147 95085 66181 95113
rect 66209 95085 66243 95113
rect 66271 95085 70019 95113
rect 70047 95085 70081 95113
rect 70109 95085 81417 95113
rect 81445 95085 81479 95113
rect 81507 95085 81541 95113
rect 81569 95085 81603 95113
rect 81631 95085 85379 95113
rect 85407 95085 85441 95113
rect 85469 95085 96777 95113
rect 96805 95085 96839 95113
rect 96867 95085 96901 95113
rect 96929 95085 96963 95113
rect 96991 95085 112137 95113
rect 112165 95085 112199 95113
rect 112227 95085 112261 95113
rect 112289 95085 112323 95113
rect 112351 95085 127497 95113
rect 127525 95085 127559 95113
rect 127587 95085 127621 95113
rect 127649 95085 127683 95113
rect 127711 95085 142857 95113
rect 142885 95085 142919 95113
rect 142947 95085 142981 95113
rect 143009 95085 143043 95113
rect 143071 95085 158217 95113
rect 158245 95085 158279 95113
rect 158307 95085 158341 95113
rect 158369 95085 158403 95113
rect 158431 95085 169939 95113
rect 169967 95085 170001 95113
rect 170029 95085 185299 95113
rect 185327 95085 185361 95113
rect 185389 95085 200659 95113
rect 200687 95085 200721 95113
rect 200749 95085 216019 95113
rect 216047 95085 216081 95113
rect 216109 95085 231379 95113
rect 231407 95085 231441 95113
rect 231469 95085 246739 95113
rect 246767 95085 246801 95113
rect 246829 95085 262099 95113
rect 262127 95085 262161 95113
rect 262189 95085 281097 95113
rect 281125 95085 281159 95113
rect 281187 95085 281221 95113
rect 281249 95085 281283 95113
rect 281311 95085 296457 95113
rect 296485 95085 296519 95113
rect 296547 95085 296581 95113
rect 296609 95085 296643 95113
rect 296671 95085 298728 95113
rect 298756 95085 298790 95113
rect 298818 95085 298852 95113
rect 298880 95085 298914 95113
rect 298942 95085 298990 95113
rect -958 95051 298990 95085
rect -958 95023 -910 95051
rect -882 95023 -848 95051
rect -820 95023 -786 95051
rect -758 95023 -724 95051
rect -696 95023 4617 95051
rect 4645 95023 4679 95051
rect 4707 95023 4741 95051
rect 4769 95023 4803 95051
rect 4831 95023 19977 95051
rect 20005 95023 20039 95051
rect 20067 95023 20101 95051
rect 20129 95023 20163 95051
rect 20191 95023 23939 95051
rect 23967 95023 24001 95051
rect 24029 95023 35337 95051
rect 35365 95023 35399 95051
rect 35427 95023 35461 95051
rect 35489 95023 35523 95051
rect 35551 95023 39299 95051
rect 39327 95023 39361 95051
rect 39389 95023 50697 95051
rect 50725 95023 50759 95051
rect 50787 95023 50821 95051
rect 50849 95023 50883 95051
rect 50911 95023 54659 95051
rect 54687 95023 54721 95051
rect 54749 95023 66057 95051
rect 66085 95023 66119 95051
rect 66147 95023 66181 95051
rect 66209 95023 66243 95051
rect 66271 95023 70019 95051
rect 70047 95023 70081 95051
rect 70109 95023 81417 95051
rect 81445 95023 81479 95051
rect 81507 95023 81541 95051
rect 81569 95023 81603 95051
rect 81631 95023 85379 95051
rect 85407 95023 85441 95051
rect 85469 95023 96777 95051
rect 96805 95023 96839 95051
rect 96867 95023 96901 95051
rect 96929 95023 96963 95051
rect 96991 95023 112137 95051
rect 112165 95023 112199 95051
rect 112227 95023 112261 95051
rect 112289 95023 112323 95051
rect 112351 95023 127497 95051
rect 127525 95023 127559 95051
rect 127587 95023 127621 95051
rect 127649 95023 127683 95051
rect 127711 95023 142857 95051
rect 142885 95023 142919 95051
rect 142947 95023 142981 95051
rect 143009 95023 143043 95051
rect 143071 95023 158217 95051
rect 158245 95023 158279 95051
rect 158307 95023 158341 95051
rect 158369 95023 158403 95051
rect 158431 95023 169939 95051
rect 169967 95023 170001 95051
rect 170029 95023 185299 95051
rect 185327 95023 185361 95051
rect 185389 95023 200659 95051
rect 200687 95023 200721 95051
rect 200749 95023 216019 95051
rect 216047 95023 216081 95051
rect 216109 95023 231379 95051
rect 231407 95023 231441 95051
rect 231469 95023 246739 95051
rect 246767 95023 246801 95051
rect 246829 95023 262099 95051
rect 262127 95023 262161 95051
rect 262189 95023 281097 95051
rect 281125 95023 281159 95051
rect 281187 95023 281221 95051
rect 281249 95023 281283 95051
rect 281311 95023 296457 95051
rect 296485 95023 296519 95051
rect 296547 95023 296581 95051
rect 296609 95023 296643 95051
rect 296671 95023 298728 95051
rect 298756 95023 298790 95051
rect 298818 95023 298852 95051
rect 298880 95023 298914 95051
rect 298942 95023 298990 95051
rect -958 94989 298990 95023
rect -958 94961 -910 94989
rect -882 94961 -848 94989
rect -820 94961 -786 94989
rect -758 94961 -724 94989
rect -696 94961 4617 94989
rect 4645 94961 4679 94989
rect 4707 94961 4741 94989
rect 4769 94961 4803 94989
rect 4831 94961 19977 94989
rect 20005 94961 20039 94989
rect 20067 94961 20101 94989
rect 20129 94961 20163 94989
rect 20191 94961 23939 94989
rect 23967 94961 24001 94989
rect 24029 94961 35337 94989
rect 35365 94961 35399 94989
rect 35427 94961 35461 94989
rect 35489 94961 35523 94989
rect 35551 94961 39299 94989
rect 39327 94961 39361 94989
rect 39389 94961 50697 94989
rect 50725 94961 50759 94989
rect 50787 94961 50821 94989
rect 50849 94961 50883 94989
rect 50911 94961 54659 94989
rect 54687 94961 54721 94989
rect 54749 94961 66057 94989
rect 66085 94961 66119 94989
rect 66147 94961 66181 94989
rect 66209 94961 66243 94989
rect 66271 94961 70019 94989
rect 70047 94961 70081 94989
rect 70109 94961 81417 94989
rect 81445 94961 81479 94989
rect 81507 94961 81541 94989
rect 81569 94961 81603 94989
rect 81631 94961 85379 94989
rect 85407 94961 85441 94989
rect 85469 94961 96777 94989
rect 96805 94961 96839 94989
rect 96867 94961 96901 94989
rect 96929 94961 96963 94989
rect 96991 94961 112137 94989
rect 112165 94961 112199 94989
rect 112227 94961 112261 94989
rect 112289 94961 112323 94989
rect 112351 94961 127497 94989
rect 127525 94961 127559 94989
rect 127587 94961 127621 94989
rect 127649 94961 127683 94989
rect 127711 94961 142857 94989
rect 142885 94961 142919 94989
rect 142947 94961 142981 94989
rect 143009 94961 143043 94989
rect 143071 94961 158217 94989
rect 158245 94961 158279 94989
rect 158307 94961 158341 94989
rect 158369 94961 158403 94989
rect 158431 94961 169939 94989
rect 169967 94961 170001 94989
rect 170029 94961 185299 94989
rect 185327 94961 185361 94989
rect 185389 94961 200659 94989
rect 200687 94961 200721 94989
rect 200749 94961 216019 94989
rect 216047 94961 216081 94989
rect 216109 94961 231379 94989
rect 231407 94961 231441 94989
rect 231469 94961 246739 94989
rect 246767 94961 246801 94989
rect 246829 94961 262099 94989
rect 262127 94961 262161 94989
rect 262189 94961 281097 94989
rect 281125 94961 281159 94989
rect 281187 94961 281221 94989
rect 281249 94961 281283 94989
rect 281311 94961 296457 94989
rect 296485 94961 296519 94989
rect 296547 94961 296581 94989
rect 296609 94961 296643 94989
rect 296671 94961 298728 94989
rect 298756 94961 298790 94989
rect 298818 94961 298852 94989
rect 298880 94961 298914 94989
rect 298942 94961 298990 94989
rect -958 94913 298990 94961
rect -958 92175 298990 92223
rect -958 92147 -430 92175
rect -402 92147 -368 92175
rect -340 92147 -306 92175
rect -278 92147 -244 92175
rect -216 92147 2757 92175
rect 2785 92147 2819 92175
rect 2847 92147 2881 92175
rect 2909 92147 2943 92175
rect 2971 92147 16259 92175
rect 16287 92147 16321 92175
rect 16349 92147 18117 92175
rect 18145 92147 18179 92175
rect 18207 92147 18241 92175
rect 18269 92147 18303 92175
rect 18331 92147 31619 92175
rect 31647 92147 31681 92175
rect 31709 92147 33477 92175
rect 33505 92147 33539 92175
rect 33567 92147 33601 92175
rect 33629 92147 33663 92175
rect 33691 92147 46979 92175
rect 47007 92147 47041 92175
rect 47069 92147 48837 92175
rect 48865 92147 48899 92175
rect 48927 92147 48961 92175
rect 48989 92147 49023 92175
rect 49051 92147 62339 92175
rect 62367 92147 62401 92175
rect 62429 92147 64197 92175
rect 64225 92147 64259 92175
rect 64287 92147 64321 92175
rect 64349 92147 64383 92175
rect 64411 92147 77699 92175
rect 77727 92147 77761 92175
rect 77789 92147 79557 92175
rect 79585 92147 79619 92175
rect 79647 92147 79681 92175
rect 79709 92147 79743 92175
rect 79771 92147 93059 92175
rect 93087 92147 93121 92175
rect 93149 92147 94917 92175
rect 94945 92147 94979 92175
rect 95007 92147 95041 92175
rect 95069 92147 95103 92175
rect 95131 92147 110277 92175
rect 110305 92147 110339 92175
rect 110367 92147 110401 92175
rect 110429 92147 110463 92175
rect 110491 92147 125637 92175
rect 125665 92147 125699 92175
rect 125727 92147 125761 92175
rect 125789 92147 125823 92175
rect 125851 92147 140997 92175
rect 141025 92147 141059 92175
rect 141087 92147 141121 92175
rect 141149 92147 141183 92175
rect 141211 92147 156357 92175
rect 156385 92147 156419 92175
rect 156447 92147 156481 92175
rect 156509 92147 156543 92175
rect 156571 92147 162259 92175
rect 162287 92147 162321 92175
rect 162349 92147 177619 92175
rect 177647 92147 177681 92175
rect 177709 92147 192979 92175
rect 193007 92147 193041 92175
rect 193069 92147 208339 92175
rect 208367 92147 208401 92175
rect 208429 92147 223699 92175
rect 223727 92147 223761 92175
rect 223789 92147 239059 92175
rect 239087 92147 239121 92175
rect 239149 92147 254419 92175
rect 254447 92147 254481 92175
rect 254509 92147 269779 92175
rect 269807 92147 269841 92175
rect 269869 92147 279237 92175
rect 279265 92147 279299 92175
rect 279327 92147 279361 92175
rect 279389 92147 279423 92175
rect 279451 92147 294597 92175
rect 294625 92147 294659 92175
rect 294687 92147 294721 92175
rect 294749 92147 294783 92175
rect 294811 92147 298248 92175
rect 298276 92147 298310 92175
rect 298338 92147 298372 92175
rect 298400 92147 298434 92175
rect 298462 92147 298990 92175
rect -958 92113 298990 92147
rect -958 92085 -430 92113
rect -402 92085 -368 92113
rect -340 92085 -306 92113
rect -278 92085 -244 92113
rect -216 92085 2757 92113
rect 2785 92085 2819 92113
rect 2847 92085 2881 92113
rect 2909 92085 2943 92113
rect 2971 92085 16259 92113
rect 16287 92085 16321 92113
rect 16349 92085 18117 92113
rect 18145 92085 18179 92113
rect 18207 92085 18241 92113
rect 18269 92085 18303 92113
rect 18331 92085 31619 92113
rect 31647 92085 31681 92113
rect 31709 92085 33477 92113
rect 33505 92085 33539 92113
rect 33567 92085 33601 92113
rect 33629 92085 33663 92113
rect 33691 92085 46979 92113
rect 47007 92085 47041 92113
rect 47069 92085 48837 92113
rect 48865 92085 48899 92113
rect 48927 92085 48961 92113
rect 48989 92085 49023 92113
rect 49051 92085 62339 92113
rect 62367 92085 62401 92113
rect 62429 92085 64197 92113
rect 64225 92085 64259 92113
rect 64287 92085 64321 92113
rect 64349 92085 64383 92113
rect 64411 92085 77699 92113
rect 77727 92085 77761 92113
rect 77789 92085 79557 92113
rect 79585 92085 79619 92113
rect 79647 92085 79681 92113
rect 79709 92085 79743 92113
rect 79771 92085 93059 92113
rect 93087 92085 93121 92113
rect 93149 92085 94917 92113
rect 94945 92085 94979 92113
rect 95007 92085 95041 92113
rect 95069 92085 95103 92113
rect 95131 92085 110277 92113
rect 110305 92085 110339 92113
rect 110367 92085 110401 92113
rect 110429 92085 110463 92113
rect 110491 92085 125637 92113
rect 125665 92085 125699 92113
rect 125727 92085 125761 92113
rect 125789 92085 125823 92113
rect 125851 92085 140997 92113
rect 141025 92085 141059 92113
rect 141087 92085 141121 92113
rect 141149 92085 141183 92113
rect 141211 92085 156357 92113
rect 156385 92085 156419 92113
rect 156447 92085 156481 92113
rect 156509 92085 156543 92113
rect 156571 92085 162259 92113
rect 162287 92085 162321 92113
rect 162349 92085 177619 92113
rect 177647 92085 177681 92113
rect 177709 92085 192979 92113
rect 193007 92085 193041 92113
rect 193069 92085 208339 92113
rect 208367 92085 208401 92113
rect 208429 92085 223699 92113
rect 223727 92085 223761 92113
rect 223789 92085 239059 92113
rect 239087 92085 239121 92113
rect 239149 92085 254419 92113
rect 254447 92085 254481 92113
rect 254509 92085 269779 92113
rect 269807 92085 269841 92113
rect 269869 92085 279237 92113
rect 279265 92085 279299 92113
rect 279327 92085 279361 92113
rect 279389 92085 279423 92113
rect 279451 92085 294597 92113
rect 294625 92085 294659 92113
rect 294687 92085 294721 92113
rect 294749 92085 294783 92113
rect 294811 92085 298248 92113
rect 298276 92085 298310 92113
rect 298338 92085 298372 92113
rect 298400 92085 298434 92113
rect 298462 92085 298990 92113
rect -958 92051 298990 92085
rect -958 92023 -430 92051
rect -402 92023 -368 92051
rect -340 92023 -306 92051
rect -278 92023 -244 92051
rect -216 92023 2757 92051
rect 2785 92023 2819 92051
rect 2847 92023 2881 92051
rect 2909 92023 2943 92051
rect 2971 92023 16259 92051
rect 16287 92023 16321 92051
rect 16349 92023 18117 92051
rect 18145 92023 18179 92051
rect 18207 92023 18241 92051
rect 18269 92023 18303 92051
rect 18331 92023 31619 92051
rect 31647 92023 31681 92051
rect 31709 92023 33477 92051
rect 33505 92023 33539 92051
rect 33567 92023 33601 92051
rect 33629 92023 33663 92051
rect 33691 92023 46979 92051
rect 47007 92023 47041 92051
rect 47069 92023 48837 92051
rect 48865 92023 48899 92051
rect 48927 92023 48961 92051
rect 48989 92023 49023 92051
rect 49051 92023 62339 92051
rect 62367 92023 62401 92051
rect 62429 92023 64197 92051
rect 64225 92023 64259 92051
rect 64287 92023 64321 92051
rect 64349 92023 64383 92051
rect 64411 92023 77699 92051
rect 77727 92023 77761 92051
rect 77789 92023 79557 92051
rect 79585 92023 79619 92051
rect 79647 92023 79681 92051
rect 79709 92023 79743 92051
rect 79771 92023 93059 92051
rect 93087 92023 93121 92051
rect 93149 92023 94917 92051
rect 94945 92023 94979 92051
rect 95007 92023 95041 92051
rect 95069 92023 95103 92051
rect 95131 92023 110277 92051
rect 110305 92023 110339 92051
rect 110367 92023 110401 92051
rect 110429 92023 110463 92051
rect 110491 92023 125637 92051
rect 125665 92023 125699 92051
rect 125727 92023 125761 92051
rect 125789 92023 125823 92051
rect 125851 92023 140997 92051
rect 141025 92023 141059 92051
rect 141087 92023 141121 92051
rect 141149 92023 141183 92051
rect 141211 92023 156357 92051
rect 156385 92023 156419 92051
rect 156447 92023 156481 92051
rect 156509 92023 156543 92051
rect 156571 92023 162259 92051
rect 162287 92023 162321 92051
rect 162349 92023 177619 92051
rect 177647 92023 177681 92051
rect 177709 92023 192979 92051
rect 193007 92023 193041 92051
rect 193069 92023 208339 92051
rect 208367 92023 208401 92051
rect 208429 92023 223699 92051
rect 223727 92023 223761 92051
rect 223789 92023 239059 92051
rect 239087 92023 239121 92051
rect 239149 92023 254419 92051
rect 254447 92023 254481 92051
rect 254509 92023 269779 92051
rect 269807 92023 269841 92051
rect 269869 92023 279237 92051
rect 279265 92023 279299 92051
rect 279327 92023 279361 92051
rect 279389 92023 279423 92051
rect 279451 92023 294597 92051
rect 294625 92023 294659 92051
rect 294687 92023 294721 92051
rect 294749 92023 294783 92051
rect 294811 92023 298248 92051
rect 298276 92023 298310 92051
rect 298338 92023 298372 92051
rect 298400 92023 298434 92051
rect 298462 92023 298990 92051
rect -958 91989 298990 92023
rect -958 91961 -430 91989
rect -402 91961 -368 91989
rect -340 91961 -306 91989
rect -278 91961 -244 91989
rect -216 91961 2757 91989
rect 2785 91961 2819 91989
rect 2847 91961 2881 91989
rect 2909 91961 2943 91989
rect 2971 91961 16259 91989
rect 16287 91961 16321 91989
rect 16349 91961 18117 91989
rect 18145 91961 18179 91989
rect 18207 91961 18241 91989
rect 18269 91961 18303 91989
rect 18331 91961 31619 91989
rect 31647 91961 31681 91989
rect 31709 91961 33477 91989
rect 33505 91961 33539 91989
rect 33567 91961 33601 91989
rect 33629 91961 33663 91989
rect 33691 91961 46979 91989
rect 47007 91961 47041 91989
rect 47069 91961 48837 91989
rect 48865 91961 48899 91989
rect 48927 91961 48961 91989
rect 48989 91961 49023 91989
rect 49051 91961 62339 91989
rect 62367 91961 62401 91989
rect 62429 91961 64197 91989
rect 64225 91961 64259 91989
rect 64287 91961 64321 91989
rect 64349 91961 64383 91989
rect 64411 91961 77699 91989
rect 77727 91961 77761 91989
rect 77789 91961 79557 91989
rect 79585 91961 79619 91989
rect 79647 91961 79681 91989
rect 79709 91961 79743 91989
rect 79771 91961 93059 91989
rect 93087 91961 93121 91989
rect 93149 91961 94917 91989
rect 94945 91961 94979 91989
rect 95007 91961 95041 91989
rect 95069 91961 95103 91989
rect 95131 91961 110277 91989
rect 110305 91961 110339 91989
rect 110367 91961 110401 91989
rect 110429 91961 110463 91989
rect 110491 91961 125637 91989
rect 125665 91961 125699 91989
rect 125727 91961 125761 91989
rect 125789 91961 125823 91989
rect 125851 91961 140997 91989
rect 141025 91961 141059 91989
rect 141087 91961 141121 91989
rect 141149 91961 141183 91989
rect 141211 91961 156357 91989
rect 156385 91961 156419 91989
rect 156447 91961 156481 91989
rect 156509 91961 156543 91989
rect 156571 91961 162259 91989
rect 162287 91961 162321 91989
rect 162349 91961 177619 91989
rect 177647 91961 177681 91989
rect 177709 91961 192979 91989
rect 193007 91961 193041 91989
rect 193069 91961 208339 91989
rect 208367 91961 208401 91989
rect 208429 91961 223699 91989
rect 223727 91961 223761 91989
rect 223789 91961 239059 91989
rect 239087 91961 239121 91989
rect 239149 91961 254419 91989
rect 254447 91961 254481 91989
rect 254509 91961 269779 91989
rect 269807 91961 269841 91989
rect 269869 91961 279237 91989
rect 279265 91961 279299 91989
rect 279327 91961 279361 91989
rect 279389 91961 279423 91989
rect 279451 91961 294597 91989
rect 294625 91961 294659 91989
rect 294687 91961 294721 91989
rect 294749 91961 294783 91989
rect 294811 91961 298248 91989
rect 298276 91961 298310 91989
rect 298338 91961 298372 91989
rect 298400 91961 298434 91989
rect 298462 91961 298990 91989
rect -958 91913 298990 91961
rect -958 86175 298990 86223
rect -958 86147 -910 86175
rect -882 86147 -848 86175
rect -820 86147 -786 86175
rect -758 86147 -724 86175
rect -696 86147 4617 86175
rect 4645 86147 4679 86175
rect 4707 86147 4741 86175
rect 4769 86147 4803 86175
rect 4831 86147 19977 86175
rect 20005 86147 20039 86175
rect 20067 86147 20101 86175
rect 20129 86147 20163 86175
rect 20191 86147 23939 86175
rect 23967 86147 24001 86175
rect 24029 86147 39299 86175
rect 39327 86147 39361 86175
rect 39389 86147 54659 86175
rect 54687 86147 54721 86175
rect 54749 86147 70019 86175
rect 70047 86147 70081 86175
rect 70109 86147 81417 86175
rect 81445 86147 81479 86175
rect 81507 86147 81541 86175
rect 81569 86147 81603 86175
rect 81631 86147 85379 86175
rect 85407 86147 85441 86175
rect 85469 86147 96777 86175
rect 96805 86147 96839 86175
rect 96867 86147 96901 86175
rect 96929 86147 96963 86175
rect 96991 86147 112137 86175
rect 112165 86147 112199 86175
rect 112227 86147 112261 86175
rect 112289 86147 112323 86175
rect 112351 86147 127497 86175
rect 127525 86147 127559 86175
rect 127587 86147 127621 86175
rect 127649 86147 127683 86175
rect 127711 86147 142857 86175
rect 142885 86147 142919 86175
rect 142947 86147 142981 86175
rect 143009 86147 143043 86175
rect 143071 86147 158217 86175
rect 158245 86147 158279 86175
rect 158307 86147 158341 86175
rect 158369 86147 158403 86175
rect 158431 86147 169939 86175
rect 169967 86147 170001 86175
rect 170029 86147 185299 86175
rect 185327 86147 185361 86175
rect 185389 86147 200659 86175
rect 200687 86147 200721 86175
rect 200749 86147 216019 86175
rect 216047 86147 216081 86175
rect 216109 86147 231379 86175
rect 231407 86147 231441 86175
rect 231469 86147 246739 86175
rect 246767 86147 246801 86175
rect 246829 86147 262099 86175
rect 262127 86147 262161 86175
rect 262189 86147 281097 86175
rect 281125 86147 281159 86175
rect 281187 86147 281221 86175
rect 281249 86147 281283 86175
rect 281311 86147 296457 86175
rect 296485 86147 296519 86175
rect 296547 86147 296581 86175
rect 296609 86147 296643 86175
rect 296671 86147 298728 86175
rect 298756 86147 298790 86175
rect 298818 86147 298852 86175
rect 298880 86147 298914 86175
rect 298942 86147 298990 86175
rect -958 86113 298990 86147
rect -958 86085 -910 86113
rect -882 86085 -848 86113
rect -820 86085 -786 86113
rect -758 86085 -724 86113
rect -696 86085 4617 86113
rect 4645 86085 4679 86113
rect 4707 86085 4741 86113
rect 4769 86085 4803 86113
rect 4831 86085 19977 86113
rect 20005 86085 20039 86113
rect 20067 86085 20101 86113
rect 20129 86085 20163 86113
rect 20191 86085 23939 86113
rect 23967 86085 24001 86113
rect 24029 86085 39299 86113
rect 39327 86085 39361 86113
rect 39389 86085 54659 86113
rect 54687 86085 54721 86113
rect 54749 86085 70019 86113
rect 70047 86085 70081 86113
rect 70109 86085 81417 86113
rect 81445 86085 81479 86113
rect 81507 86085 81541 86113
rect 81569 86085 81603 86113
rect 81631 86085 85379 86113
rect 85407 86085 85441 86113
rect 85469 86085 96777 86113
rect 96805 86085 96839 86113
rect 96867 86085 96901 86113
rect 96929 86085 96963 86113
rect 96991 86085 112137 86113
rect 112165 86085 112199 86113
rect 112227 86085 112261 86113
rect 112289 86085 112323 86113
rect 112351 86085 127497 86113
rect 127525 86085 127559 86113
rect 127587 86085 127621 86113
rect 127649 86085 127683 86113
rect 127711 86085 142857 86113
rect 142885 86085 142919 86113
rect 142947 86085 142981 86113
rect 143009 86085 143043 86113
rect 143071 86085 158217 86113
rect 158245 86085 158279 86113
rect 158307 86085 158341 86113
rect 158369 86085 158403 86113
rect 158431 86085 169939 86113
rect 169967 86085 170001 86113
rect 170029 86085 185299 86113
rect 185327 86085 185361 86113
rect 185389 86085 200659 86113
rect 200687 86085 200721 86113
rect 200749 86085 216019 86113
rect 216047 86085 216081 86113
rect 216109 86085 231379 86113
rect 231407 86085 231441 86113
rect 231469 86085 246739 86113
rect 246767 86085 246801 86113
rect 246829 86085 262099 86113
rect 262127 86085 262161 86113
rect 262189 86085 281097 86113
rect 281125 86085 281159 86113
rect 281187 86085 281221 86113
rect 281249 86085 281283 86113
rect 281311 86085 296457 86113
rect 296485 86085 296519 86113
rect 296547 86085 296581 86113
rect 296609 86085 296643 86113
rect 296671 86085 298728 86113
rect 298756 86085 298790 86113
rect 298818 86085 298852 86113
rect 298880 86085 298914 86113
rect 298942 86085 298990 86113
rect -958 86051 298990 86085
rect -958 86023 -910 86051
rect -882 86023 -848 86051
rect -820 86023 -786 86051
rect -758 86023 -724 86051
rect -696 86023 4617 86051
rect 4645 86023 4679 86051
rect 4707 86023 4741 86051
rect 4769 86023 4803 86051
rect 4831 86023 19977 86051
rect 20005 86023 20039 86051
rect 20067 86023 20101 86051
rect 20129 86023 20163 86051
rect 20191 86023 23939 86051
rect 23967 86023 24001 86051
rect 24029 86023 39299 86051
rect 39327 86023 39361 86051
rect 39389 86023 54659 86051
rect 54687 86023 54721 86051
rect 54749 86023 70019 86051
rect 70047 86023 70081 86051
rect 70109 86023 81417 86051
rect 81445 86023 81479 86051
rect 81507 86023 81541 86051
rect 81569 86023 81603 86051
rect 81631 86023 85379 86051
rect 85407 86023 85441 86051
rect 85469 86023 96777 86051
rect 96805 86023 96839 86051
rect 96867 86023 96901 86051
rect 96929 86023 96963 86051
rect 96991 86023 112137 86051
rect 112165 86023 112199 86051
rect 112227 86023 112261 86051
rect 112289 86023 112323 86051
rect 112351 86023 127497 86051
rect 127525 86023 127559 86051
rect 127587 86023 127621 86051
rect 127649 86023 127683 86051
rect 127711 86023 142857 86051
rect 142885 86023 142919 86051
rect 142947 86023 142981 86051
rect 143009 86023 143043 86051
rect 143071 86023 158217 86051
rect 158245 86023 158279 86051
rect 158307 86023 158341 86051
rect 158369 86023 158403 86051
rect 158431 86023 169939 86051
rect 169967 86023 170001 86051
rect 170029 86023 185299 86051
rect 185327 86023 185361 86051
rect 185389 86023 200659 86051
rect 200687 86023 200721 86051
rect 200749 86023 216019 86051
rect 216047 86023 216081 86051
rect 216109 86023 231379 86051
rect 231407 86023 231441 86051
rect 231469 86023 246739 86051
rect 246767 86023 246801 86051
rect 246829 86023 262099 86051
rect 262127 86023 262161 86051
rect 262189 86023 281097 86051
rect 281125 86023 281159 86051
rect 281187 86023 281221 86051
rect 281249 86023 281283 86051
rect 281311 86023 296457 86051
rect 296485 86023 296519 86051
rect 296547 86023 296581 86051
rect 296609 86023 296643 86051
rect 296671 86023 298728 86051
rect 298756 86023 298790 86051
rect 298818 86023 298852 86051
rect 298880 86023 298914 86051
rect 298942 86023 298990 86051
rect -958 85989 298990 86023
rect -958 85961 -910 85989
rect -882 85961 -848 85989
rect -820 85961 -786 85989
rect -758 85961 -724 85989
rect -696 85961 4617 85989
rect 4645 85961 4679 85989
rect 4707 85961 4741 85989
rect 4769 85961 4803 85989
rect 4831 85961 19977 85989
rect 20005 85961 20039 85989
rect 20067 85961 20101 85989
rect 20129 85961 20163 85989
rect 20191 85961 23939 85989
rect 23967 85961 24001 85989
rect 24029 85961 39299 85989
rect 39327 85961 39361 85989
rect 39389 85961 54659 85989
rect 54687 85961 54721 85989
rect 54749 85961 70019 85989
rect 70047 85961 70081 85989
rect 70109 85961 81417 85989
rect 81445 85961 81479 85989
rect 81507 85961 81541 85989
rect 81569 85961 81603 85989
rect 81631 85961 85379 85989
rect 85407 85961 85441 85989
rect 85469 85961 96777 85989
rect 96805 85961 96839 85989
rect 96867 85961 96901 85989
rect 96929 85961 96963 85989
rect 96991 85961 112137 85989
rect 112165 85961 112199 85989
rect 112227 85961 112261 85989
rect 112289 85961 112323 85989
rect 112351 85961 127497 85989
rect 127525 85961 127559 85989
rect 127587 85961 127621 85989
rect 127649 85961 127683 85989
rect 127711 85961 142857 85989
rect 142885 85961 142919 85989
rect 142947 85961 142981 85989
rect 143009 85961 143043 85989
rect 143071 85961 158217 85989
rect 158245 85961 158279 85989
rect 158307 85961 158341 85989
rect 158369 85961 158403 85989
rect 158431 85961 169939 85989
rect 169967 85961 170001 85989
rect 170029 85961 185299 85989
rect 185327 85961 185361 85989
rect 185389 85961 200659 85989
rect 200687 85961 200721 85989
rect 200749 85961 216019 85989
rect 216047 85961 216081 85989
rect 216109 85961 231379 85989
rect 231407 85961 231441 85989
rect 231469 85961 246739 85989
rect 246767 85961 246801 85989
rect 246829 85961 262099 85989
rect 262127 85961 262161 85989
rect 262189 85961 281097 85989
rect 281125 85961 281159 85989
rect 281187 85961 281221 85989
rect 281249 85961 281283 85989
rect 281311 85961 296457 85989
rect 296485 85961 296519 85989
rect 296547 85961 296581 85989
rect 296609 85961 296643 85989
rect 296671 85961 298728 85989
rect 298756 85961 298790 85989
rect 298818 85961 298852 85989
rect 298880 85961 298914 85989
rect 298942 85961 298990 85989
rect -958 85913 298990 85961
rect -958 83175 298990 83223
rect -958 83147 -430 83175
rect -402 83147 -368 83175
rect -340 83147 -306 83175
rect -278 83147 -244 83175
rect -216 83147 2757 83175
rect 2785 83147 2819 83175
rect 2847 83147 2881 83175
rect 2909 83147 2943 83175
rect 2971 83147 16259 83175
rect 16287 83147 16321 83175
rect 16349 83147 18117 83175
rect 18145 83147 18179 83175
rect 18207 83147 18241 83175
rect 18269 83147 18303 83175
rect 18331 83147 31619 83175
rect 31647 83147 31681 83175
rect 31709 83147 46979 83175
rect 47007 83147 47041 83175
rect 47069 83147 62339 83175
rect 62367 83147 62401 83175
rect 62429 83147 77699 83175
rect 77727 83147 77761 83175
rect 77789 83147 79557 83175
rect 79585 83147 79619 83175
rect 79647 83147 79681 83175
rect 79709 83147 79743 83175
rect 79771 83147 93059 83175
rect 93087 83147 93121 83175
rect 93149 83147 94917 83175
rect 94945 83147 94979 83175
rect 95007 83147 95041 83175
rect 95069 83147 95103 83175
rect 95131 83147 110277 83175
rect 110305 83147 110339 83175
rect 110367 83147 110401 83175
rect 110429 83147 110463 83175
rect 110491 83147 125637 83175
rect 125665 83147 125699 83175
rect 125727 83147 125761 83175
rect 125789 83147 125823 83175
rect 125851 83147 140997 83175
rect 141025 83147 141059 83175
rect 141087 83147 141121 83175
rect 141149 83147 141183 83175
rect 141211 83147 156357 83175
rect 156385 83147 156419 83175
rect 156447 83147 156481 83175
rect 156509 83147 156543 83175
rect 156571 83147 162259 83175
rect 162287 83147 162321 83175
rect 162349 83147 177619 83175
rect 177647 83147 177681 83175
rect 177709 83147 192979 83175
rect 193007 83147 193041 83175
rect 193069 83147 208339 83175
rect 208367 83147 208401 83175
rect 208429 83147 223699 83175
rect 223727 83147 223761 83175
rect 223789 83147 239059 83175
rect 239087 83147 239121 83175
rect 239149 83147 254419 83175
rect 254447 83147 254481 83175
rect 254509 83147 269779 83175
rect 269807 83147 269841 83175
rect 269869 83147 279237 83175
rect 279265 83147 279299 83175
rect 279327 83147 279361 83175
rect 279389 83147 279423 83175
rect 279451 83147 294597 83175
rect 294625 83147 294659 83175
rect 294687 83147 294721 83175
rect 294749 83147 294783 83175
rect 294811 83147 298248 83175
rect 298276 83147 298310 83175
rect 298338 83147 298372 83175
rect 298400 83147 298434 83175
rect 298462 83147 298990 83175
rect -958 83113 298990 83147
rect -958 83085 -430 83113
rect -402 83085 -368 83113
rect -340 83085 -306 83113
rect -278 83085 -244 83113
rect -216 83085 2757 83113
rect 2785 83085 2819 83113
rect 2847 83085 2881 83113
rect 2909 83085 2943 83113
rect 2971 83085 16259 83113
rect 16287 83085 16321 83113
rect 16349 83085 18117 83113
rect 18145 83085 18179 83113
rect 18207 83085 18241 83113
rect 18269 83085 18303 83113
rect 18331 83085 31619 83113
rect 31647 83085 31681 83113
rect 31709 83085 46979 83113
rect 47007 83085 47041 83113
rect 47069 83085 62339 83113
rect 62367 83085 62401 83113
rect 62429 83085 77699 83113
rect 77727 83085 77761 83113
rect 77789 83085 79557 83113
rect 79585 83085 79619 83113
rect 79647 83085 79681 83113
rect 79709 83085 79743 83113
rect 79771 83085 93059 83113
rect 93087 83085 93121 83113
rect 93149 83085 94917 83113
rect 94945 83085 94979 83113
rect 95007 83085 95041 83113
rect 95069 83085 95103 83113
rect 95131 83085 110277 83113
rect 110305 83085 110339 83113
rect 110367 83085 110401 83113
rect 110429 83085 110463 83113
rect 110491 83085 125637 83113
rect 125665 83085 125699 83113
rect 125727 83085 125761 83113
rect 125789 83085 125823 83113
rect 125851 83085 140997 83113
rect 141025 83085 141059 83113
rect 141087 83085 141121 83113
rect 141149 83085 141183 83113
rect 141211 83085 156357 83113
rect 156385 83085 156419 83113
rect 156447 83085 156481 83113
rect 156509 83085 156543 83113
rect 156571 83085 162259 83113
rect 162287 83085 162321 83113
rect 162349 83085 177619 83113
rect 177647 83085 177681 83113
rect 177709 83085 192979 83113
rect 193007 83085 193041 83113
rect 193069 83085 208339 83113
rect 208367 83085 208401 83113
rect 208429 83085 223699 83113
rect 223727 83085 223761 83113
rect 223789 83085 239059 83113
rect 239087 83085 239121 83113
rect 239149 83085 254419 83113
rect 254447 83085 254481 83113
rect 254509 83085 269779 83113
rect 269807 83085 269841 83113
rect 269869 83085 279237 83113
rect 279265 83085 279299 83113
rect 279327 83085 279361 83113
rect 279389 83085 279423 83113
rect 279451 83085 294597 83113
rect 294625 83085 294659 83113
rect 294687 83085 294721 83113
rect 294749 83085 294783 83113
rect 294811 83085 298248 83113
rect 298276 83085 298310 83113
rect 298338 83085 298372 83113
rect 298400 83085 298434 83113
rect 298462 83085 298990 83113
rect -958 83051 298990 83085
rect -958 83023 -430 83051
rect -402 83023 -368 83051
rect -340 83023 -306 83051
rect -278 83023 -244 83051
rect -216 83023 2757 83051
rect 2785 83023 2819 83051
rect 2847 83023 2881 83051
rect 2909 83023 2943 83051
rect 2971 83023 16259 83051
rect 16287 83023 16321 83051
rect 16349 83023 18117 83051
rect 18145 83023 18179 83051
rect 18207 83023 18241 83051
rect 18269 83023 18303 83051
rect 18331 83023 31619 83051
rect 31647 83023 31681 83051
rect 31709 83023 46979 83051
rect 47007 83023 47041 83051
rect 47069 83023 62339 83051
rect 62367 83023 62401 83051
rect 62429 83023 77699 83051
rect 77727 83023 77761 83051
rect 77789 83023 79557 83051
rect 79585 83023 79619 83051
rect 79647 83023 79681 83051
rect 79709 83023 79743 83051
rect 79771 83023 93059 83051
rect 93087 83023 93121 83051
rect 93149 83023 94917 83051
rect 94945 83023 94979 83051
rect 95007 83023 95041 83051
rect 95069 83023 95103 83051
rect 95131 83023 110277 83051
rect 110305 83023 110339 83051
rect 110367 83023 110401 83051
rect 110429 83023 110463 83051
rect 110491 83023 125637 83051
rect 125665 83023 125699 83051
rect 125727 83023 125761 83051
rect 125789 83023 125823 83051
rect 125851 83023 140997 83051
rect 141025 83023 141059 83051
rect 141087 83023 141121 83051
rect 141149 83023 141183 83051
rect 141211 83023 156357 83051
rect 156385 83023 156419 83051
rect 156447 83023 156481 83051
rect 156509 83023 156543 83051
rect 156571 83023 162259 83051
rect 162287 83023 162321 83051
rect 162349 83023 177619 83051
rect 177647 83023 177681 83051
rect 177709 83023 192979 83051
rect 193007 83023 193041 83051
rect 193069 83023 208339 83051
rect 208367 83023 208401 83051
rect 208429 83023 223699 83051
rect 223727 83023 223761 83051
rect 223789 83023 239059 83051
rect 239087 83023 239121 83051
rect 239149 83023 254419 83051
rect 254447 83023 254481 83051
rect 254509 83023 269779 83051
rect 269807 83023 269841 83051
rect 269869 83023 279237 83051
rect 279265 83023 279299 83051
rect 279327 83023 279361 83051
rect 279389 83023 279423 83051
rect 279451 83023 294597 83051
rect 294625 83023 294659 83051
rect 294687 83023 294721 83051
rect 294749 83023 294783 83051
rect 294811 83023 298248 83051
rect 298276 83023 298310 83051
rect 298338 83023 298372 83051
rect 298400 83023 298434 83051
rect 298462 83023 298990 83051
rect -958 82989 298990 83023
rect -958 82961 -430 82989
rect -402 82961 -368 82989
rect -340 82961 -306 82989
rect -278 82961 -244 82989
rect -216 82961 2757 82989
rect 2785 82961 2819 82989
rect 2847 82961 2881 82989
rect 2909 82961 2943 82989
rect 2971 82961 16259 82989
rect 16287 82961 16321 82989
rect 16349 82961 18117 82989
rect 18145 82961 18179 82989
rect 18207 82961 18241 82989
rect 18269 82961 18303 82989
rect 18331 82961 31619 82989
rect 31647 82961 31681 82989
rect 31709 82961 46979 82989
rect 47007 82961 47041 82989
rect 47069 82961 62339 82989
rect 62367 82961 62401 82989
rect 62429 82961 77699 82989
rect 77727 82961 77761 82989
rect 77789 82961 79557 82989
rect 79585 82961 79619 82989
rect 79647 82961 79681 82989
rect 79709 82961 79743 82989
rect 79771 82961 93059 82989
rect 93087 82961 93121 82989
rect 93149 82961 94917 82989
rect 94945 82961 94979 82989
rect 95007 82961 95041 82989
rect 95069 82961 95103 82989
rect 95131 82961 110277 82989
rect 110305 82961 110339 82989
rect 110367 82961 110401 82989
rect 110429 82961 110463 82989
rect 110491 82961 125637 82989
rect 125665 82961 125699 82989
rect 125727 82961 125761 82989
rect 125789 82961 125823 82989
rect 125851 82961 140997 82989
rect 141025 82961 141059 82989
rect 141087 82961 141121 82989
rect 141149 82961 141183 82989
rect 141211 82961 156357 82989
rect 156385 82961 156419 82989
rect 156447 82961 156481 82989
rect 156509 82961 156543 82989
rect 156571 82961 162259 82989
rect 162287 82961 162321 82989
rect 162349 82961 177619 82989
rect 177647 82961 177681 82989
rect 177709 82961 192979 82989
rect 193007 82961 193041 82989
rect 193069 82961 208339 82989
rect 208367 82961 208401 82989
rect 208429 82961 223699 82989
rect 223727 82961 223761 82989
rect 223789 82961 239059 82989
rect 239087 82961 239121 82989
rect 239149 82961 254419 82989
rect 254447 82961 254481 82989
rect 254509 82961 269779 82989
rect 269807 82961 269841 82989
rect 269869 82961 279237 82989
rect 279265 82961 279299 82989
rect 279327 82961 279361 82989
rect 279389 82961 279423 82989
rect 279451 82961 294597 82989
rect 294625 82961 294659 82989
rect 294687 82961 294721 82989
rect 294749 82961 294783 82989
rect 294811 82961 298248 82989
rect 298276 82961 298310 82989
rect 298338 82961 298372 82989
rect 298400 82961 298434 82989
rect 298462 82961 298990 82989
rect -958 82913 298990 82961
rect -958 77175 298990 77223
rect -958 77147 -910 77175
rect -882 77147 -848 77175
rect -820 77147 -786 77175
rect -758 77147 -724 77175
rect -696 77147 4617 77175
rect 4645 77147 4679 77175
rect 4707 77147 4741 77175
rect 4769 77147 4803 77175
rect 4831 77147 19977 77175
rect 20005 77147 20039 77175
rect 20067 77147 20101 77175
rect 20129 77147 20163 77175
rect 20191 77147 23939 77175
rect 23967 77147 24001 77175
rect 24029 77147 39299 77175
rect 39327 77147 39361 77175
rect 39389 77147 54659 77175
rect 54687 77147 54721 77175
rect 54749 77147 70019 77175
rect 70047 77147 70081 77175
rect 70109 77147 81417 77175
rect 81445 77147 81479 77175
rect 81507 77147 81541 77175
rect 81569 77147 81603 77175
rect 81631 77147 85379 77175
rect 85407 77147 85441 77175
rect 85469 77147 96777 77175
rect 96805 77147 96839 77175
rect 96867 77147 96901 77175
rect 96929 77147 96963 77175
rect 96991 77147 112137 77175
rect 112165 77147 112199 77175
rect 112227 77147 112261 77175
rect 112289 77147 112323 77175
rect 112351 77147 127497 77175
rect 127525 77147 127559 77175
rect 127587 77147 127621 77175
rect 127649 77147 127683 77175
rect 127711 77147 142857 77175
rect 142885 77147 142919 77175
rect 142947 77147 142981 77175
rect 143009 77147 143043 77175
rect 143071 77147 158217 77175
rect 158245 77147 158279 77175
rect 158307 77147 158341 77175
rect 158369 77147 158403 77175
rect 158431 77147 169939 77175
rect 169967 77147 170001 77175
rect 170029 77147 185299 77175
rect 185327 77147 185361 77175
rect 185389 77147 200659 77175
rect 200687 77147 200721 77175
rect 200749 77147 216019 77175
rect 216047 77147 216081 77175
rect 216109 77147 231379 77175
rect 231407 77147 231441 77175
rect 231469 77147 246739 77175
rect 246767 77147 246801 77175
rect 246829 77147 262099 77175
rect 262127 77147 262161 77175
rect 262189 77147 281097 77175
rect 281125 77147 281159 77175
rect 281187 77147 281221 77175
rect 281249 77147 281283 77175
rect 281311 77147 296457 77175
rect 296485 77147 296519 77175
rect 296547 77147 296581 77175
rect 296609 77147 296643 77175
rect 296671 77147 298728 77175
rect 298756 77147 298790 77175
rect 298818 77147 298852 77175
rect 298880 77147 298914 77175
rect 298942 77147 298990 77175
rect -958 77113 298990 77147
rect -958 77085 -910 77113
rect -882 77085 -848 77113
rect -820 77085 -786 77113
rect -758 77085 -724 77113
rect -696 77085 4617 77113
rect 4645 77085 4679 77113
rect 4707 77085 4741 77113
rect 4769 77085 4803 77113
rect 4831 77085 19977 77113
rect 20005 77085 20039 77113
rect 20067 77085 20101 77113
rect 20129 77085 20163 77113
rect 20191 77085 23939 77113
rect 23967 77085 24001 77113
rect 24029 77085 39299 77113
rect 39327 77085 39361 77113
rect 39389 77085 54659 77113
rect 54687 77085 54721 77113
rect 54749 77085 70019 77113
rect 70047 77085 70081 77113
rect 70109 77085 81417 77113
rect 81445 77085 81479 77113
rect 81507 77085 81541 77113
rect 81569 77085 81603 77113
rect 81631 77085 85379 77113
rect 85407 77085 85441 77113
rect 85469 77085 96777 77113
rect 96805 77085 96839 77113
rect 96867 77085 96901 77113
rect 96929 77085 96963 77113
rect 96991 77085 112137 77113
rect 112165 77085 112199 77113
rect 112227 77085 112261 77113
rect 112289 77085 112323 77113
rect 112351 77085 127497 77113
rect 127525 77085 127559 77113
rect 127587 77085 127621 77113
rect 127649 77085 127683 77113
rect 127711 77085 142857 77113
rect 142885 77085 142919 77113
rect 142947 77085 142981 77113
rect 143009 77085 143043 77113
rect 143071 77085 158217 77113
rect 158245 77085 158279 77113
rect 158307 77085 158341 77113
rect 158369 77085 158403 77113
rect 158431 77085 169939 77113
rect 169967 77085 170001 77113
rect 170029 77085 185299 77113
rect 185327 77085 185361 77113
rect 185389 77085 200659 77113
rect 200687 77085 200721 77113
rect 200749 77085 216019 77113
rect 216047 77085 216081 77113
rect 216109 77085 231379 77113
rect 231407 77085 231441 77113
rect 231469 77085 246739 77113
rect 246767 77085 246801 77113
rect 246829 77085 262099 77113
rect 262127 77085 262161 77113
rect 262189 77085 281097 77113
rect 281125 77085 281159 77113
rect 281187 77085 281221 77113
rect 281249 77085 281283 77113
rect 281311 77085 296457 77113
rect 296485 77085 296519 77113
rect 296547 77085 296581 77113
rect 296609 77085 296643 77113
rect 296671 77085 298728 77113
rect 298756 77085 298790 77113
rect 298818 77085 298852 77113
rect 298880 77085 298914 77113
rect 298942 77085 298990 77113
rect -958 77051 298990 77085
rect -958 77023 -910 77051
rect -882 77023 -848 77051
rect -820 77023 -786 77051
rect -758 77023 -724 77051
rect -696 77023 4617 77051
rect 4645 77023 4679 77051
rect 4707 77023 4741 77051
rect 4769 77023 4803 77051
rect 4831 77023 19977 77051
rect 20005 77023 20039 77051
rect 20067 77023 20101 77051
rect 20129 77023 20163 77051
rect 20191 77023 23939 77051
rect 23967 77023 24001 77051
rect 24029 77023 39299 77051
rect 39327 77023 39361 77051
rect 39389 77023 54659 77051
rect 54687 77023 54721 77051
rect 54749 77023 70019 77051
rect 70047 77023 70081 77051
rect 70109 77023 81417 77051
rect 81445 77023 81479 77051
rect 81507 77023 81541 77051
rect 81569 77023 81603 77051
rect 81631 77023 85379 77051
rect 85407 77023 85441 77051
rect 85469 77023 96777 77051
rect 96805 77023 96839 77051
rect 96867 77023 96901 77051
rect 96929 77023 96963 77051
rect 96991 77023 112137 77051
rect 112165 77023 112199 77051
rect 112227 77023 112261 77051
rect 112289 77023 112323 77051
rect 112351 77023 127497 77051
rect 127525 77023 127559 77051
rect 127587 77023 127621 77051
rect 127649 77023 127683 77051
rect 127711 77023 142857 77051
rect 142885 77023 142919 77051
rect 142947 77023 142981 77051
rect 143009 77023 143043 77051
rect 143071 77023 158217 77051
rect 158245 77023 158279 77051
rect 158307 77023 158341 77051
rect 158369 77023 158403 77051
rect 158431 77023 169939 77051
rect 169967 77023 170001 77051
rect 170029 77023 185299 77051
rect 185327 77023 185361 77051
rect 185389 77023 200659 77051
rect 200687 77023 200721 77051
rect 200749 77023 216019 77051
rect 216047 77023 216081 77051
rect 216109 77023 231379 77051
rect 231407 77023 231441 77051
rect 231469 77023 246739 77051
rect 246767 77023 246801 77051
rect 246829 77023 262099 77051
rect 262127 77023 262161 77051
rect 262189 77023 281097 77051
rect 281125 77023 281159 77051
rect 281187 77023 281221 77051
rect 281249 77023 281283 77051
rect 281311 77023 296457 77051
rect 296485 77023 296519 77051
rect 296547 77023 296581 77051
rect 296609 77023 296643 77051
rect 296671 77023 298728 77051
rect 298756 77023 298790 77051
rect 298818 77023 298852 77051
rect 298880 77023 298914 77051
rect 298942 77023 298990 77051
rect -958 76989 298990 77023
rect -958 76961 -910 76989
rect -882 76961 -848 76989
rect -820 76961 -786 76989
rect -758 76961 -724 76989
rect -696 76961 4617 76989
rect 4645 76961 4679 76989
rect 4707 76961 4741 76989
rect 4769 76961 4803 76989
rect 4831 76961 19977 76989
rect 20005 76961 20039 76989
rect 20067 76961 20101 76989
rect 20129 76961 20163 76989
rect 20191 76961 23939 76989
rect 23967 76961 24001 76989
rect 24029 76961 39299 76989
rect 39327 76961 39361 76989
rect 39389 76961 54659 76989
rect 54687 76961 54721 76989
rect 54749 76961 70019 76989
rect 70047 76961 70081 76989
rect 70109 76961 81417 76989
rect 81445 76961 81479 76989
rect 81507 76961 81541 76989
rect 81569 76961 81603 76989
rect 81631 76961 85379 76989
rect 85407 76961 85441 76989
rect 85469 76961 96777 76989
rect 96805 76961 96839 76989
rect 96867 76961 96901 76989
rect 96929 76961 96963 76989
rect 96991 76961 112137 76989
rect 112165 76961 112199 76989
rect 112227 76961 112261 76989
rect 112289 76961 112323 76989
rect 112351 76961 127497 76989
rect 127525 76961 127559 76989
rect 127587 76961 127621 76989
rect 127649 76961 127683 76989
rect 127711 76961 142857 76989
rect 142885 76961 142919 76989
rect 142947 76961 142981 76989
rect 143009 76961 143043 76989
rect 143071 76961 158217 76989
rect 158245 76961 158279 76989
rect 158307 76961 158341 76989
rect 158369 76961 158403 76989
rect 158431 76961 169939 76989
rect 169967 76961 170001 76989
rect 170029 76961 185299 76989
rect 185327 76961 185361 76989
rect 185389 76961 200659 76989
rect 200687 76961 200721 76989
rect 200749 76961 216019 76989
rect 216047 76961 216081 76989
rect 216109 76961 231379 76989
rect 231407 76961 231441 76989
rect 231469 76961 246739 76989
rect 246767 76961 246801 76989
rect 246829 76961 262099 76989
rect 262127 76961 262161 76989
rect 262189 76961 281097 76989
rect 281125 76961 281159 76989
rect 281187 76961 281221 76989
rect 281249 76961 281283 76989
rect 281311 76961 296457 76989
rect 296485 76961 296519 76989
rect 296547 76961 296581 76989
rect 296609 76961 296643 76989
rect 296671 76961 298728 76989
rect 298756 76961 298790 76989
rect 298818 76961 298852 76989
rect 298880 76961 298914 76989
rect 298942 76961 298990 76989
rect -958 76913 298990 76961
rect -958 74175 298990 74223
rect -958 74147 -430 74175
rect -402 74147 -368 74175
rect -340 74147 -306 74175
rect -278 74147 -244 74175
rect -216 74147 2757 74175
rect 2785 74147 2819 74175
rect 2847 74147 2881 74175
rect 2909 74147 2943 74175
rect 2971 74147 18117 74175
rect 18145 74147 18179 74175
rect 18207 74147 18241 74175
rect 18269 74147 18303 74175
rect 18331 74147 33477 74175
rect 33505 74147 33539 74175
rect 33567 74147 33601 74175
rect 33629 74147 33663 74175
rect 33691 74147 48837 74175
rect 48865 74147 48899 74175
rect 48927 74147 48961 74175
rect 48989 74147 49023 74175
rect 49051 74147 64197 74175
rect 64225 74147 64259 74175
rect 64287 74147 64321 74175
rect 64349 74147 64383 74175
rect 64411 74147 79557 74175
rect 79585 74147 79619 74175
rect 79647 74147 79681 74175
rect 79709 74147 79743 74175
rect 79771 74147 94917 74175
rect 94945 74147 94979 74175
rect 95007 74147 95041 74175
rect 95069 74147 95103 74175
rect 95131 74147 110277 74175
rect 110305 74147 110339 74175
rect 110367 74147 110401 74175
rect 110429 74147 110463 74175
rect 110491 74147 125637 74175
rect 125665 74147 125699 74175
rect 125727 74147 125761 74175
rect 125789 74147 125823 74175
rect 125851 74147 140997 74175
rect 141025 74147 141059 74175
rect 141087 74147 141121 74175
rect 141149 74147 141183 74175
rect 141211 74147 156357 74175
rect 156385 74147 156419 74175
rect 156447 74147 156481 74175
rect 156509 74147 156543 74175
rect 156571 74147 162259 74175
rect 162287 74147 162321 74175
rect 162349 74147 177619 74175
rect 177647 74147 177681 74175
rect 177709 74147 192979 74175
rect 193007 74147 193041 74175
rect 193069 74147 208339 74175
rect 208367 74147 208401 74175
rect 208429 74147 223699 74175
rect 223727 74147 223761 74175
rect 223789 74147 239059 74175
rect 239087 74147 239121 74175
rect 239149 74147 254419 74175
rect 254447 74147 254481 74175
rect 254509 74147 269779 74175
rect 269807 74147 269841 74175
rect 269869 74147 279237 74175
rect 279265 74147 279299 74175
rect 279327 74147 279361 74175
rect 279389 74147 279423 74175
rect 279451 74147 294597 74175
rect 294625 74147 294659 74175
rect 294687 74147 294721 74175
rect 294749 74147 294783 74175
rect 294811 74147 298248 74175
rect 298276 74147 298310 74175
rect 298338 74147 298372 74175
rect 298400 74147 298434 74175
rect 298462 74147 298990 74175
rect -958 74113 298990 74147
rect -958 74085 -430 74113
rect -402 74085 -368 74113
rect -340 74085 -306 74113
rect -278 74085 -244 74113
rect -216 74085 2757 74113
rect 2785 74085 2819 74113
rect 2847 74085 2881 74113
rect 2909 74085 2943 74113
rect 2971 74085 18117 74113
rect 18145 74085 18179 74113
rect 18207 74085 18241 74113
rect 18269 74085 18303 74113
rect 18331 74085 33477 74113
rect 33505 74085 33539 74113
rect 33567 74085 33601 74113
rect 33629 74085 33663 74113
rect 33691 74085 48837 74113
rect 48865 74085 48899 74113
rect 48927 74085 48961 74113
rect 48989 74085 49023 74113
rect 49051 74085 64197 74113
rect 64225 74085 64259 74113
rect 64287 74085 64321 74113
rect 64349 74085 64383 74113
rect 64411 74085 79557 74113
rect 79585 74085 79619 74113
rect 79647 74085 79681 74113
rect 79709 74085 79743 74113
rect 79771 74085 94917 74113
rect 94945 74085 94979 74113
rect 95007 74085 95041 74113
rect 95069 74085 95103 74113
rect 95131 74085 110277 74113
rect 110305 74085 110339 74113
rect 110367 74085 110401 74113
rect 110429 74085 110463 74113
rect 110491 74085 125637 74113
rect 125665 74085 125699 74113
rect 125727 74085 125761 74113
rect 125789 74085 125823 74113
rect 125851 74085 140997 74113
rect 141025 74085 141059 74113
rect 141087 74085 141121 74113
rect 141149 74085 141183 74113
rect 141211 74085 156357 74113
rect 156385 74085 156419 74113
rect 156447 74085 156481 74113
rect 156509 74085 156543 74113
rect 156571 74085 162259 74113
rect 162287 74085 162321 74113
rect 162349 74085 177619 74113
rect 177647 74085 177681 74113
rect 177709 74085 192979 74113
rect 193007 74085 193041 74113
rect 193069 74085 208339 74113
rect 208367 74085 208401 74113
rect 208429 74085 223699 74113
rect 223727 74085 223761 74113
rect 223789 74085 239059 74113
rect 239087 74085 239121 74113
rect 239149 74085 254419 74113
rect 254447 74085 254481 74113
rect 254509 74085 269779 74113
rect 269807 74085 269841 74113
rect 269869 74085 279237 74113
rect 279265 74085 279299 74113
rect 279327 74085 279361 74113
rect 279389 74085 279423 74113
rect 279451 74085 294597 74113
rect 294625 74085 294659 74113
rect 294687 74085 294721 74113
rect 294749 74085 294783 74113
rect 294811 74085 298248 74113
rect 298276 74085 298310 74113
rect 298338 74085 298372 74113
rect 298400 74085 298434 74113
rect 298462 74085 298990 74113
rect -958 74051 298990 74085
rect -958 74023 -430 74051
rect -402 74023 -368 74051
rect -340 74023 -306 74051
rect -278 74023 -244 74051
rect -216 74023 2757 74051
rect 2785 74023 2819 74051
rect 2847 74023 2881 74051
rect 2909 74023 2943 74051
rect 2971 74023 18117 74051
rect 18145 74023 18179 74051
rect 18207 74023 18241 74051
rect 18269 74023 18303 74051
rect 18331 74023 33477 74051
rect 33505 74023 33539 74051
rect 33567 74023 33601 74051
rect 33629 74023 33663 74051
rect 33691 74023 48837 74051
rect 48865 74023 48899 74051
rect 48927 74023 48961 74051
rect 48989 74023 49023 74051
rect 49051 74023 64197 74051
rect 64225 74023 64259 74051
rect 64287 74023 64321 74051
rect 64349 74023 64383 74051
rect 64411 74023 79557 74051
rect 79585 74023 79619 74051
rect 79647 74023 79681 74051
rect 79709 74023 79743 74051
rect 79771 74023 94917 74051
rect 94945 74023 94979 74051
rect 95007 74023 95041 74051
rect 95069 74023 95103 74051
rect 95131 74023 110277 74051
rect 110305 74023 110339 74051
rect 110367 74023 110401 74051
rect 110429 74023 110463 74051
rect 110491 74023 125637 74051
rect 125665 74023 125699 74051
rect 125727 74023 125761 74051
rect 125789 74023 125823 74051
rect 125851 74023 140997 74051
rect 141025 74023 141059 74051
rect 141087 74023 141121 74051
rect 141149 74023 141183 74051
rect 141211 74023 156357 74051
rect 156385 74023 156419 74051
rect 156447 74023 156481 74051
rect 156509 74023 156543 74051
rect 156571 74023 162259 74051
rect 162287 74023 162321 74051
rect 162349 74023 177619 74051
rect 177647 74023 177681 74051
rect 177709 74023 192979 74051
rect 193007 74023 193041 74051
rect 193069 74023 208339 74051
rect 208367 74023 208401 74051
rect 208429 74023 223699 74051
rect 223727 74023 223761 74051
rect 223789 74023 239059 74051
rect 239087 74023 239121 74051
rect 239149 74023 254419 74051
rect 254447 74023 254481 74051
rect 254509 74023 269779 74051
rect 269807 74023 269841 74051
rect 269869 74023 279237 74051
rect 279265 74023 279299 74051
rect 279327 74023 279361 74051
rect 279389 74023 279423 74051
rect 279451 74023 294597 74051
rect 294625 74023 294659 74051
rect 294687 74023 294721 74051
rect 294749 74023 294783 74051
rect 294811 74023 298248 74051
rect 298276 74023 298310 74051
rect 298338 74023 298372 74051
rect 298400 74023 298434 74051
rect 298462 74023 298990 74051
rect -958 73989 298990 74023
rect -958 73961 -430 73989
rect -402 73961 -368 73989
rect -340 73961 -306 73989
rect -278 73961 -244 73989
rect -216 73961 2757 73989
rect 2785 73961 2819 73989
rect 2847 73961 2881 73989
rect 2909 73961 2943 73989
rect 2971 73961 18117 73989
rect 18145 73961 18179 73989
rect 18207 73961 18241 73989
rect 18269 73961 18303 73989
rect 18331 73961 33477 73989
rect 33505 73961 33539 73989
rect 33567 73961 33601 73989
rect 33629 73961 33663 73989
rect 33691 73961 48837 73989
rect 48865 73961 48899 73989
rect 48927 73961 48961 73989
rect 48989 73961 49023 73989
rect 49051 73961 64197 73989
rect 64225 73961 64259 73989
rect 64287 73961 64321 73989
rect 64349 73961 64383 73989
rect 64411 73961 79557 73989
rect 79585 73961 79619 73989
rect 79647 73961 79681 73989
rect 79709 73961 79743 73989
rect 79771 73961 94917 73989
rect 94945 73961 94979 73989
rect 95007 73961 95041 73989
rect 95069 73961 95103 73989
rect 95131 73961 110277 73989
rect 110305 73961 110339 73989
rect 110367 73961 110401 73989
rect 110429 73961 110463 73989
rect 110491 73961 125637 73989
rect 125665 73961 125699 73989
rect 125727 73961 125761 73989
rect 125789 73961 125823 73989
rect 125851 73961 140997 73989
rect 141025 73961 141059 73989
rect 141087 73961 141121 73989
rect 141149 73961 141183 73989
rect 141211 73961 156357 73989
rect 156385 73961 156419 73989
rect 156447 73961 156481 73989
rect 156509 73961 156543 73989
rect 156571 73961 162259 73989
rect 162287 73961 162321 73989
rect 162349 73961 177619 73989
rect 177647 73961 177681 73989
rect 177709 73961 192979 73989
rect 193007 73961 193041 73989
rect 193069 73961 208339 73989
rect 208367 73961 208401 73989
rect 208429 73961 223699 73989
rect 223727 73961 223761 73989
rect 223789 73961 239059 73989
rect 239087 73961 239121 73989
rect 239149 73961 254419 73989
rect 254447 73961 254481 73989
rect 254509 73961 269779 73989
rect 269807 73961 269841 73989
rect 269869 73961 279237 73989
rect 279265 73961 279299 73989
rect 279327 73961 279361 73989
rect 279389 73961 279423 73989
rect 279451 73961 294597 73989
rect 294625 73961 294659 73989
rect 294687 73961 294721 73989
rect 294749 73961 294783 73989
rect 294811 73961 298248 73989
rect 298276 73961 298310 73989
rect 298338 73961 298372 73989
rect 298400 73961 298434 73989
rect 298462 73961 298990 73989
rect -958 73913 298990 73961
rect -958 68175 298990 68223
rect -958 68147 -910 68175
rect -882 68147 -848 68175
rect -820 68147 -786 68175
rect -758 68147 -724 68175
rect -696 68147 4617 68175
rect 4645 68147 4679 68175
rect 4707 68147 4741 68175
rect 4769 68147 4803 68175
rect 4831 68147 19977 68175
rect 20005 68147 20039 68175
rect 20067 68147 20101 68175
rect 20129 68147 20163 68175
rect 20191 68147 35337 68175
rect 35365 68147 35399 68175
rect 35427 68147 35461 68175
rect 35489 68147 35523 68175
rect 35551 68147 50697 68175
rect 50725 68147 50759 68175
rect 50787 68147 50821 68175
rect 50849 68147 50883 68175
rect 50911 68147 66057 68175
rect 66085 68147 66119 68175
rect 66147 68147 66181 68175
rect 66209 68147 66243 68175
rect 66271 68147 81417 68175
rect 81445 68147 81479 68175
rect 81507 68147 81541 68175
rect 81569 68147 81603 68175
rect 81631 68147 96777 68175
rect 96805 68147 96839 68175
rect 96867 68147 96901 68175
rect 96929 68147 96963 68175
rect 96991 68147 112137 68175
rect 112165 68147 112199 68175
rect 112227 68147 112261 68175
rect 112289 68147 112323 68175
rect 112351 68147 127497 68175
rect 127525 68147 127559 68175
rect 127587 68147 127621 68175
rect 127649 68147 127683 68175
rect 127711 68147 142857 68175
rect 142885 68147 142919 68175
rect 142947 68147 142981 68175
rect 143009 68147 143043 68175
rect 143071 68147 158217 68175
rect 158245 68147 158279 68175
rect 158307 68147 158341 68175
rect 158369 68147 158403 68175
rect 158431 68147 169939 68175
rect 169967 68147 170001 68175
rect 170029 68147 185299 68175
rect 185327 68147 185361 68175
rect 185389 68147 200659 68175
rect 200687 68147 200721 68175
rect 200749 68147 216019 68175
rect 216047 68147 216081 68175
rect 216109 68147 231379 68175
rect 231407 68147 231441 68175
rect 231469 68147 246739 68175
rect 246767 68147 246801 68175
rect 246829 68147 262099 68175
rect 262127 68147 262161 68175
rect 262189 68147 281097 68175
rect 281125 68147 281159 68175
rect 281187 68147 281221 68175
rect 281249 68147 281283 68175
rect 281311 68147 296457 68175
rect 296485 68147 296519 68175
rect 296547 68147 296581 68175
rect 296609 68147 296643 68175
rect 296671 68147 298728 68175
rect 298756 68147 298790 68175
rect 298818 68147 298852 68175
rect 298880 68147 298914 68175
rect 298942 68147 298990 68175
rect -958 68113 298990 68147
rect -958 68085 -910 68113
rect -882 68085 -848 68113
rect -820 68085 -786 68113
rect -758 68085 -724 68113
rect -696 68085 4617 68113
rect 4645 68085 4679 68113
rect 4707 68085 4741 68113
rect 4769 68085 4803 68113
rect 4831 68085 19977 68113
rect 20005 68085 20039 68113
rect 20067 68085 20101 68113
rect 20129 68085 20163 68113
rect 20191 68085 35337 68113
rect 35365 68085 35399 68113
rect 35427 68085 35461 68113
rect 35489 68085 35523 68113
rect 35551 68085 50697 68113
rect 50725 68085 50759 68113
rect 50787 68085 50821 68113
rect 50849 68085 50883 68113
rect 50911 68085 66057 68113
rect 66085 68085 66119 68113
rect 66147 68085 66181 68113
rect 66209 68085 66243 68113
rect 66271 68085 81417 68113
rect 81445 68085 81479 68113
rect 81507 68085 81541 68113
rect 81569 68085 81603 68113
rect 81631 68085 96777 68113
rect 96805 68085 96839 68113
rect 96867 68085 96901 68113
rect 96929 68085 96963 68113
rect 96991 68085 112137 68113
rect 112165 68085 112199 68113
rect 112227 68085 112261 68113
rect 112289 68085 112323 68113
rect 112351 68085 127497 68113
rect 127525 68085 127559 68113
rect 127587 68085 127621 68113
rect 127649 68085 127683 68113
rect 127711 68085 142857 68113
rect 142885 68085 142919 68113
rect 142947 68085 142981 68113
rect 143009 68085 143043 68113
rect 143071 68085 158217 68113
rect 158245 68085 158279 68113
rect 158307 68085 158341 68113
rect 158369 68085 158403 68113
rect 158431 68085 169939 68113
rect 169967 68085 170001 68113
rect 170029 68085 185299 68113
rect 185327 68085 185361 68113
rect 185389 68085 200659 68113
rect 200687 68085 200721 68113
rect 200749 68085 216019 68113
rect 216047 68085 216081 68113
rect 216109 68085 231379 68113
rect 231407 68085 231441 68113
rect 231469 68085 246739 68113
rect 246767 68085 246801 68113
rect 246829 68085 262099 68113
rect 262127 68085 262161 68113
rect 262189 68085 281097 68113
rect 281125 68085 281159 68113
rect 281187 68085 281221 68113
rect 281249 68085 281283 68113
rect 281311 68085 296457 68113
rect 296485 68085 296519 68113
rect 296547 68085 296581 68113
rect 296609 68085 296643 68113
rect 296671 68085 298728 68113
rect 298756 68085 298790 68113
rect 298818 68085 298852 68113
rect 298880 68085 298914 68113
rect 298942 68085 298990 68113
rect -958 68051 298990 68085
rect -958 68023 -910 68051
rect -882 68023 -848 68051
rect -820 68023 -786 68051
rect -758 68023 -724 68051
rect -696 68023 4617 68051
rect 4645 68023 4679 68051
rect 4707 68023 4741 68051
rect 4769 68023 4803 68051
rect 4831 68023 19977 68051
rect 20005 68023 20039 68051
rect 20067 68023 20101 68051
rect 20129 68023 20163 68051
rect 20191 68023 35337 68051
rect 35365 68023 35399 68051
rect 35427 68023 35461 68051
rect 35489 68023 35523 68051
rect 35551 68023 50697 68051
rect 50725 68023 50759 68051
rect 50787 68023 50821 68051
rect 50849 68023 50883 68051
rect 50911 68023 66057 68051
rect 66085 68023 66119 68051
rect 66147 68023 66181 68051
rect 66209 68023 66243 68051
rect 66271 68023 81417 68051
rect 81445 68023 81479 68051
rect 81507 68023 81541 68051
rect 81569 68023 81603 68051
rect 81631 68023 96777 68051
rect 96805 68023 96839 68051
rect 96867 68023 96901 68051
rect 96929 68023 96963 68051
rect 96991 68023 112137 68051
rect 112165 68023 112199 68051
rect 112227 68023 112261 68051
rect 112289 68023 112323 68051
rect 112351 68023 127497 68051
rect 127525 68023 127559 68051
rect 127587 68023 127621 68051
rect 127649 68023 127683 68051
rect 127711 68023 142857 68051
rect 142885 68023 142919 68051
rect 142947 68023 142981 68051
rect 143009 68023 143043 68051
rect 143071 68023 158217 68051
rect 158245 68023 158279 68051
rect 158307 68023 158341 68051
rect 158369 68023 158403 68051
rect 158431 68023 169939 68051
rect 169967 68023 170001 68051
rect 170029 68023 185299 68051
rect 185327 68023 185361 68051
rect 185389 68023 200659 68051
rect 200687 68023 200721 68051
rect 200749 68023 216019 68051
rect 216047 68023 216081 68051
rect 216109 68023 231379 68051
rect 231407 68023 231441 68051
rect 231469 68023 246739 68051
rect 246767 68023 246801 68051
rect 246829 68023 262099 68051
rect 262127 68023 262161 68051
rect 262189 68023 281097 68051
rect 281125 68023 281159 68051
rect 281187 68023 281221 68051
rect 281249 68023 281283 68051
rect 281311 68023 296457 68051
rect 296485 68023 296519 68051
rect 296547 68023 296581 68051
rect 296609 68023 296643 68051
rect 296671 68023 298728 68051
rect 298756 68023 298790 68051
rect 298818 68023 298852 68051
rect 298880 68023 298914 68051
rect 298942 68023 298990 68051
rect -958 67989 298990 68023
rect -958 67961 -910 67989
rect -882 67961 -848 67989
rect -820 67961 -786 67989
rect -758 67961 -724 67989
rect -696 67961 4617 67989
rect 4645 67961 4679 67989
rect 4707 67961 4741 67989
rect 4769 67961 4803 67989
rect 4831 67961 19977 67989
rect 20005 67961 20039 67989
rect 20067 67961 20101 67989
rect 20129 67961 20163 67989
rect 20191 67961 35337 67989
rect 35365 67961 35399 67989
rect 35427 67961 35461 67989
rect 35489 67961 35523 67989
rect 35551 67961 50697 67989
rect 50725 67961 50759 67989
rect 50787 67961 50821 67989
rect 50849 67961 50883 67989
rect 50911 67961 66057 67989
rect 66085 67961 66119 67989
rect 66147 67961 66181 67989
rect 66209 67961 66243 67989
rect 66271 67961 81417 67989
rect 81445 67961 81479 67989
rect 81507 67961 81541 67989
rect 81569 67961 81603 67989
rect 81631 67961 96777 67989
rect 96805 67961 96839 67989
rect 96867 67961 96901 67989
rect 96929 67961 96963 67989
rect 96991 67961 112137 67989
rect 112165 67961 112199 67989
rect 112227 67961 112261 67989
rect 112289 67961 112323 67989
rect 112351 67961 127497 67989
rect 127525 67961 127559 67989
rect 127587 67961 127621 67989
rect 127649 67961 127683 67989
rect 127711 67961 142857 67989
rect 142885 67961 142919 67989
rect 142947 67961 142981 67989
rect 143009 67961 143043 67989
rect 143071 67961 158217 67989
rect 158245 67961 158279 67989
rect 158307 67961 158341 67989
rect 158369 67961 158403 67989
rect 158431 67961 169939 67989
rect 169967 67961 170001 67989
rect 170029 67961 185299 67989
rect 185327 67961 185361 67989
rect 185389 67961 200659 67989
rect 200687 67961 200721 67989
rect 200749 67961 216019 67989
rect 216047 67961 216081 67989
rect 216109 67961 231379 67989
rect 231407 67961 231441 67989
rect 231469 67961 246739 67989
rect 246767 67961 246801 67989
rect 246829 67961 262099 67989
rect 262127 67961 262161 67989
rect 262189 67961 281097 67989
rect 281125 67961 281159 67989
rect 281187 67961 281221 67989
rect 281249 67961 281283 67989
rect 281311 67961 296457 67989
rect 296485 67961 296519 67989
rect 296547 67961 296581 67989
rect 296609 67961 296643 67989
rect 296671 67961 298728 67989
rect 298756 67961 298790 67989
rect 298818 67961 298852 67989
rect 298880 67961 298914 67989
rect 298942 67961 298990 67989
rect -958 67913 298990 67961
rect -958 65175 298990 65223
rect -958 65147 -430 65175
rect -402 65147 -368 65175
rect -340 65147 -306 65175
rect -278 65147 -244 65175
rect -216 65147 2757 65175
rect 2785 65147 2819 65175
rect 2847 65147 2881 65175
rect 2909 65147 2943 65175
rect 2971 65147 18117 65175
rect 18145 65147 18179 65175
rect 18207 65147 18241 65175
rect 18269 65147 18303 65175
rect 18331 65147 33477 65175
rect 33505 65147 33539 65175
rect 33567 65147 33601 65175
rect 33629 65147 33663 65175
rect 33691 65147 48837 65175
rect 48865 65147 48899 65175
rect 48927 65147 48961 65175
rect 48989 65147 49023 65175
rect 49051 65147 64197 65175
rect 64225 65147 64259 65175
rect 64287 65147 64321 65175
rect 64349 65147 64383 65175
rect 64411 65147 79557 65175
rect 79585 65147 79619 65175
rect 79647 65147 79681 65175
rect 79709 65147 79743 65175
rect 79771 65147 94917 65175
rect 94945 65147 94979 65175
rect 95007 65147 95041 65175
rect 95069 65147 95103 65175
rect 95131 65147 110277 65175
rect 110305 65147 110339 65175
rect 110367 65147 110401 65175
rect 110429 65147 110463 65175
rect 110491 65147 125637 65175
rect 125665 65147 125699 65175
rect 125727 65147 125761 65175
rect 125789 65147 125823 65175
rect 125851 65147 140997 65175
rect 141025 65147 141059 65175
rect 141087 65147 141121 65175
rect 141149 65147 141183 65175
rect 141211 65147 156357 65175
rect 156385 65147 156419 65175
rect 156447 65147 156481 65175
rect 156509 65147 156543 65175
rect 156571 65147 162259 65175
rect 162287 65147 162321 65175
rect 162349 65147 177619 65175
rect 177647 65147 177681 65175
rect 177709 65147 192979 65175
rect 193007 65147 193041 65175
rect 193069 65147 208339 65175
rect 208367 65147 208401 65175
rect 208429 65147 223699 65175
rect 223727 65147 223761 65175
rect 223789 65147 239059 65175
rect 239087 65147 239121 65175
rect 239149 65147 254419 65175
rect 254447 65147 254481 65175
rect 254509 65147 269779 65175
rect 269807 65147 269841 65175
rect 269869 65147 279237 65175
rect 279265 65147 279299 65175
rect 279327 65147 279361 65175
rect 279389 65147 279423 65175
rect 279451 65147 294597 65175
rect 294625 65147 294659 65175
rect 294687 65147 294721 65175
rect 294749 65147 294783 65175
rect 294811 65147 298248 65175
rect 298276 65147 298310 65175
rect 298338 65147 298372 65175
rect 298400 65147 298434 65175
rect 298462 65147 298990 65175
rect -958 65113 298990 65147
rect -958 65085 -430 65113
rect -402 65085 -368 65113
rect -340 65085 -306 65113
rect -278 65085 -244 65113
rect -216 65085 2757 65113
rect 2785 65085 2819 65113
rect 2847 65085 2881 65113
rect 2909 65085 2943 65113
rect 2971 65085 18117 65113
rect 18145 65085 18179 65113
rect 18207 65085 18241 65113
rect 18269 65085 18303 65113
rect 18331 65085 33477 65113
rect 33505 65085 33539 65113
rect 33567 65085 33601 65113
rect 33629 65085 33663 65113
rect 33691 65085 48837 65113
rect 48865 65085 48899 65113
rect 48927 65085 48961 65113
rect 48989 65085 49023 65113
rect 49051 65085 64197 65113
rect 64225 65085 64259 65113
rect 64287 65085 64321 65113
rect 64349 65085 64383 65113
rect 64411 65085 79557 65113
rect 79585 65085 79619 65113
rect 79647 65085 79681 65113
rect 79709 65085 79743 65113
rect 79771 65085 94917 65113
rect 94945 65085 94979 65113
rect 95007 65085 95041 65113
rect 95069 65085 95103 65113
rect 95131 65085 110277 65113
rect 110305 65085 110339 65113
rect 110367 65085 110401 65113
rect 110429 65085 110463 65113
rect 110491 65085 125637 65113
rect 125665 65085 125699 65113
rect 125727 65085 125761 65113
rect 125789 65085 125823 65113
rect 125851 65085 140997 65113
rect 141025 65085 141059 65113
rect 141087 65085 141121 65113
rect 141149 65085 141183 65113
rect 141211 65085 156357 65113
rect 156385 65085 156419 65113
rect 156447 65085 156481 65113
rect 156509 65085 156543 65113
rect 156571 65085 162259 65113
rect 162287 65085 162321 65113
rect 162349 65085 177619 65113
rect 177647 65085 177681 65113
rect 177709 65085 192979 65113
rect 193007 65085 193041 65113
rect 193069 65085 208339 65113
rect 208367 65085 208401 65113
rect 208429 65085 223699 65113
rect 223727 65085 223761 65113
rect 223789 65085 239059 65113
rect 239087 65085 239121 65113
rect 239149 65085 254419 65113
rect 254447 65085 254481 65113
rect 254509 65085 269779 65113
rect 269807 65085 269841 65113
rect 269869 65085 279237 65113
rect 279265 65085 279299 65113
rect 279327 65085 279361 65113
rect 279389 65085 279423 65113
rect 279451 65085 294597 65113
rect 294625 65085 294659 65113
rect 294687 65085 294721 65113
rect 294749 65085 294783 65113
rect 294811 65085 298248 65113
rect 298276 65085 298310 65113
rect 298338 65085 298372 65113
rect 298400 65085 298434 65113
rect 298462 65085 298990 65113
rect -958 65051 298990 65085
rect -958 65023 -430 65051
rect -402 65023 -368 65051
rect -340 65023 -306 65051
rect -278 65023 -244 65051
rect -216 65023 2757 65051
rect 2785 65023 2819 65051
rect 2847 65023 2881 65051
rect 2909 65023 2943 65051
rect 2971 65023 18117 65051
rect 18145 65023 18179 65051
rect 18207 65023 18241 65051
rect 18269 65023 18303 65051
rect 18331 65023 33477 65051
rect 33505 65023 33539 65051
rect 33567 65023 33601 65051
rect 33629 65023 33663 65051
rect 33691 65023 48837 65051
rect 48865 65023 48899 65051
rect 48927 65023 48961 65051
rect 48989 65023 49023 65051
rect 49051 65023 64197 65051
rect 64225 65023 64259 65051
rect 64287 65023 64321 65051
rect 64349 65023 64383 65051
rect 64411 65023 79557 65051
rect 79585 65023 79619 65051
rect 79647 65023 79681 65051
rect 79709 65023 79743 65051
rect 79771 65023 94917 65051
rect 94945 65023 94979 65051
rect 95007 65023 95041 65051
rect 95069 65023 95103 65051
rect 95131 65023 110277 65051
rect 110305 65023 110339 65051
rect 110367 65023 110401 65051
rect 110429 65023 110463 65051
rect 110491 65023 125637 65051
rect 125665 65023 125699 65051
rect 125727 65023 125761 65051
rect 125789 65023 125823 65051
rect 125851 65023 140997 65051
rect 141025 65023 141059 65051
rect 141087 65023 141121 65051
rect 141149 65023 141183 65051
rect 141211 65023 156357 65051
rect 156385 65023 156419 65051
rect 156447 65023 156481 65051
rect 156509 65023 156543 65051
rect 156571 65023 162259 65051
rect 162287 65023 162321 65051
rect 162349 65023 177619 65051
rect 177647 65023 177681 65051
rect 177709 65023 192979 65051
rect 193007 65023 193041 65051
rect 193069 65023 208339 65051
rect 208367 65023 208401 65051
rect 208429 65023 223699 65051
rect 223727 65023 223761 65051
rect 223789 65023 239059 65051
rect 239087 65023 239121 65051
rect 239149 65023 254419 65051
rect 254447 65023 254481 65051
rect 254509 65023 269779 65051
rect 269807 65023 269841 65051
rect 269869 65023 279237 65051
rect 279265 65023 279299 65051
rect 279327 65023 279361 65051
rect 279389 65023 279423 65051
rect 279451 65023 294597 65051
rect 294625 65023 294659 65051
rect 294687 65023 294721 65051
rect 294749 65023 294783 65051
rect 294811 65023 298248 65051
rect 298276 65023 298310 65051
rect 298338 65023 298372 65051
rect 298400 65023 298434 65051
rect 298462 65023 298990 65051
rect -958 64989 298990 65023
rect -958 64961 -430 64989
rect -402 64961 -368 64989
rect -340 64961 -306 64989
rect -278 64961 -244 64989
rect -216 64961 2757 64989
rect 2785 64961 2819 64989
rect 2847 64961 2881 64989
rect 2909 64961 2943 64989
rect 2971 64961 18117 64989
rect 18145 64961 18179 64989
rect 18207 64961 18241 64989
rect 18269 64961 18303 64989
rect 18331 64961 33477 64989
rect 33505 64961 33539 64989
rect 33567 64961 33601 64989
rect 33629 64961 33663 64989
rect 33691 64961 48837 64989
rect 48865 64961 48899 64989
rect 48927 64961 48961 64989
rect 48989 64961 49023 64989
rect 49051 64961 64197 64989
rect 64225 64961 64259 64989
rect 64287 64961 64321 64989
rect 64349 64961 64383 64989
rect 64411 64961 79557 64989
rect 79585 64961 79619 64989
rect 79647 64961 79681 64989
rect 79709 64961 79743 64989
rect 79771 64961 94917 64989
rect 94945 64961 94979 64989
rect 95007 64961 95041 64989
rect 95069 64961 95103 64989
rect 95131 64961 110277 64989
rect 110305 64961 110339 64989
rect 110367 64961 110401 64989
rect 110429 64961 110463 64989
rect 110491 64961 125637 64989
rect 125665 64961 125699 64989
rect 125727 64961 125761 64989
rect 125789 64961 125823 64989
rect 125851 64961 140997 64989
rect 141025 64961 141059 64989
rect 141087 64961 141121 64989
rect 141149 64961 141183 64989
rect 141211 64961 156357 64989
rect 156385 64961 156419 64989
rect 156447 64961 156481 64989
rect 156509 64961 156543 64989
rect 156571 64961 162259 64989
rect 162287 64961 162321 64989
rect 162349 64961 177619 64989
rect 177647 64961 177681 64989
rect 177709 64961 192979 64989
rect 193007 64961 193041 64989
rect 193069 64961 208339 64989
rect 208367 64961 208401 64989
rect 208429 64961 223699 64989
rect 223727 64961 223761 64989
rect 223789 64961 239059 64989
rect 239087 64961 239121 64989
rect 239149 64961 254419 64989
rect 254447 64961 254481 64989
rect 254509 64961 269779 64989
rect 269807 64961 269841 64989
rect 269869 64961 279237 64989
rect 279265 64961 279299 64989
rect 279327 64961 279361 64989
rect 279389 64961 279423 64989
rect 279451 64961 294597 64989
rect 294625 64961 294659 64989
rect 294687 64961 294721 64989
rect 294749 64961 294783 64989
rect 294811 64961 298248 64989
rect 298276 64961 298310 64989
rect 298338 64961 298372 64989
rect 298400 64961 298434 64989
rect 298462 64961 298990 64989
rect -958 64913 298990 64961
rect -958 59175 298990 59223
rect -958 59147 -910 59175
rect -882 59147 -848 59175
rect -820 59147 -786 59175
rect -758 59147 -724 59175
rect -696 59147 4617 59175
rect 4645 59147 4679 59175
rect 4707 59147 4741 59175
rect 4769 59147 4803 59175
rect 4831 59147 19977 59175
rect 20005 59147 20039 59175
rect 20067 59147 20101 59175
rect 20129 59147 20163 59175
rect 20191 59147 35337 59175
rect 35365 59147 35399 59175
rect 35427 59147 35461 59175
rect 35489 59147 35523 59175
rect 35551 59147 50697 59175
rect 50725 59147 50759 59175
rect 50787 59147 50821 59175
rect 50849 59147 50883 59175
rect 50911 59147 66057 59175
rect 66085 59147 66119 59175
rect 66147 59147 66181 59175
rect 66209 59147 66243 59175
rect 66271 59147 81417 59175
rect 81445 59147 81479 59175
rect 81507 59147 81541 59175
rect 81569 59147 81603 59175
rect 81631 59147 96777 59175
rect 96805 59147 96839 59175
rect 96867 59147 96901 59175
rect 96929 59147 96963 59175
rect 96991 59147 112137 59175
rect 112165 59147 112199 59175
rect 112227 59147 112261 59175
rect 112289 59147 112323 59175
rect 112351 59147 127497 59175
rect 127525 59147 127559 59175
rect 127587 59147 127621 59175
rect 127649 59147 127683 59175
rect 127711 59147 142857 59175
rect 142885 59147 142919 59175
rect 142947 59147 142981 59175
rect 143009 59147 143043 59175
rect 143071 59147 158217 59175
rect 158245 59147 158279 59175
rect 158307 59147 158341 59175
rect 158369 59147 158403 59175
rect 158431 59147 169939 59175
rect 169967 59147 170001 59175
rect 170029 59147 185299 59175
rect 185327 59147 185361 59175
rect 185389 59147 200659 59175
rect 200687 59147 200721 59175
rect 200749 59147 216019 59175
rect 216047 59147 216081 59175
rect 216109 59147 231379 59175
rect 231407 59147 231441 59175
rect 231469 59147 246739 59175
rect 246767 59147 246801 59175
rect 246829 59147 262099 59175
rect 262127 59147 262161 59175
rect 262189 59147 281097 59175
rect 281125 59147 281159 59175
rect 281187 59147 281221 59175
rect 281249 59147 281283 59175
rect 281311 59147 296457 59175
rect 296485 59147 296519 59175
rect 296547 59147 296581 59175
rect 296609 59147 296643 59175
rect 296671 59147 298728 59175
rect 298756 59147 298790 59175
rect 298818 59147 298852 59175
rect 298880 59147 298914 59175
rect 298942 59147 298990 59175
rect -958 59113 298990 59147
rect -958 59085 -910 59113
rect -882 59085 -848 59113
rect -820 59085 -786 59113
rect -758 59085 -724 59113
rect -696 59085 4617 59113
rect 4645 59085 4679 59113
rect 4707 59085 4741 59113
rect 4769 59085 4803 59113
rect 4831 59085 19977 59113
rect 20005 59085 20039 59113
rect 20067 59085 20101 59113
rect 20129 59085 20163 59113
rect 20191 59085 35337 59113
rect 35365 59085 35399 59113
rect 35427 59085 35461 59113
rect 35489 59085 35523 59113
rect 35551 59085 50697 59113
rect 50725 59085 50759 59113
rect 50787 59085 50821 59113
rect 50849 59085 50883 59113
rect 50911 59085 66057 59113
rect 66085 59085 66119 59113
rect 66147 59085 66181 59113
rect 66209 59085 66243 59113
rect 66271 59085 81417 59113
rect 81445 59085 81479 59113
rect 81507 59085 81541 59113
rect 81569 59085 81603 59113
rect 81631 59085 96777 59113
rect 96805 59085 96839 59113
rect 96867 59085 96901 59113
rect 96929 59085 96963 59113
rect 96991 59085 112137 59113
rect 112165 59085 112199 59113
rect 112227 59085 112261 59113
rect 112289 59085 112323 59113
rect 112351 59085 127497 59113
rect 127525 59085 127559 59113
rect 127587 59085 127621 59113
rect 127649 59085 127683 59113
rect 127711 59085 142857 59113
rect 142885 59085 142919 59113
rect 142947 59085 142981 59113
rect 143009 59085 143043 59113
rect 143071 59085 158217 59113
rect 158245 59085 158279 59113
rect 158307 59085 158341 59113
rect 158369 59085 158403 59113
rect 158431 59085 169939 59113
rect 169967 59085 170001 59113
rect 170029 59085 185299 59113
rect 185327 59085 185361 59113
rect 185389 59085 200659 59113
rect 200687 59085 200721 59113
rect 200749 59085 216019 59113
rect 216047 59085 216081 59113
rect 216109 59085 231379 59113
rect 231407 59085 231441 59113
rect 231469 59085 246739 59113
rect 246767 59085 246801 59113
rect 246829 59085 262099 59113
rect 262127 59085 262161 59113
rect 262189 59085 281097 59113
rect 281125 59085 281159 59113
rect 281187 59085 281221 59113
rect 281249 59085 281283 59113
rect 281311 59085 296457 59113
rect 296485 59085 296519 59113
rect 296547 59085 296581 59113
rect 296609 59085 296643 59113
rect 296671 59085 298728 59113
rect 298756 59085 298790 59113
rect 298818 59085 298852 59113
rect 298880 59085 298914 59113
rect 298942 59085 298990 59113
rect -958 59051 298990 59085
rect -958 59023 -910 59051
rect -882 59023 -848 59051
rect -820 59023 -786 59051
rect -758 59023 -724 59051
rect -696 59023 4617 59051
rect 4645 59023 4679 59051
rect 4707 59023 4741 59051
rect 4769 59023 4803 59051
rect 4831 59023 19977 59051
rect 20005 59023 20039 59051
rect 20067 59023 20101 59051
rect 20129 59023 20163 59051
rect 20191 59023 35337 59051
rect 35365 59023 35399 59051
rect 35427 59023 35461 59051
rect 35489 59023 35523 59051
rect 35551 59023 50697 59051
rect 50725 59023 50759 59051
rect 50787 59023 50821 59051
rect 50849 59023 50883 59051
rect 50911 59023 66057 59051
rect 66085 59023 66119 59051
rect 66147 59023 66181 59051
rect 66209 59023 66243 59051
rect 66271 59023 81417 59051
rect 81445 59023 81479 59051
rect 81507 59023 81541 59051
rect 81569 59023 81603 59051
rect 81631 59023 96777 59051
rect 96805 59023 96839 59051
rect 96867 59023 96901 59051
rect 96929 59023 96963 59051
rect 96991 59023 112137 59051
rect 112165 59023 112199 59051
rect 112227 59023 112261 59051
rect 112289 59023 112323 59051
rect 112351 59023 127497 59051
rect 127525 59023 127559 59051
rect 127587 59023 127621 59051
rect 127649 59023 127683 59051
rect 127711 59023 142857 59051
rect 142885 59023 142919 59051
rect 142947 59023 142981 59051
rect 143009 59023 143043 59051
rect 143071 59023 158217 59051
rect 158245 59023 158279 59051
rect 158307 59023 158341 59051
rect 158369 59023 158403 59051
rect 158431 59023 169939 59051
rect 169967 59023 170001 59051
rect 170029 59023 185299 59051
rect 185327 59023 185361 59051
rect 185389 59023 200659 59051
rect 200687 59023 200721 59051
rect 200749 59023 216019 59051
rect 216047 59023 216081 59051
rect 216109 59023 231379 59051
rect 231407 59023 231441 59051
rect 231469 59023 246739 59051
rect 246767 59023 246801 59051
rect 246829 59023 262099 59051
rect 262127 59023 262161 59051
rect 262189 59023 281097 59051
rect 281125 59023 281159 59051
rect 281187 59023 281221 59051
rect 281249 59023 281283 59051
rect 281311 59023 296457 59051
rect 296485 59023 296519 59051
rect 296547 59023 296581 59051
rect 296609 59023 296643 59051
rect 296671 59023 298728 59051
rect 298756 59023 298790 59051
rect 298818 59023 298852 59051
rect 298880 59023 298914 59051
rect 298942 59023 298990 59051
rect -958 58989 298990 59023
rect -958 58961 -910 58989
rect -882 58961 -848 58989
rect -820 58961 -786 58989
rect -758 58961 -724 58989
rect -696 58961 4617 58989
rect 4645 58961 4679 58989
rect 4707 58961 4741 58989
rect 4769 58961 4803 58989
rect 4831 58961 19977 58989
rect 20005 58961 20039 58989
rect 20067 58961 20101 58989
rect 20129 58961 20163 58989
rect 20191 58961 35337 58989
rect 35365 58961 35399 58989
rect 35427 58961 35461 58989
rect 35489 58961 35523 58989
rect 35551 58961 50697 58989
rect 50725 58961 50759 58989
rect 50787 58961 50821 58989
rect 50849 58961 50883 58989
rect 50911 58961 66057 58989
rect 66085 58961 66119 58989
rect 66147 58961 66181 58989
rect 66209 58961 66243 58989
rect 66271 58961 81417 58989
rect 81445 58961 81479 58989
rect 81507 58961 81541 58989
rect 81569 58961 81603 58989
rect 81631 58961 96777 58989
rect 96805 58961 96839 58989
rect 96867 58961 96901 58989
rect 96929 58961 96963 58989
rect 96991 58961 112137 58989
rect 112165 58961 112199 58989
rect 112227 58961 112261 58989
rect 112289 58961 112323 58989
rect 112351 58961 127497 58989
rect 127525 58961 127559 58989
rect 127587 58961 127621 58989
rect 127649 58961 127683 58989
rect 127711 58961 142857 58989
rect 142885 58961 142919 58989
rect 142947 58961 142981 58989
rect 143009 58961 143043 58989
rect 143071 58961 158217 58989
rect 158245 58961 158279 58989
rect 158307 58961 158341 58989
rect 158369 58961 158403 58989
rect 158431 58961 169939 58989
rect 169967 58961 170001 58989
rect 170029 58961 185299 58989
rect 185327 58961 185361 58989
rect 185389 58961 200659 58989
rect 200687 58961 200721 58989
rect 200749 58961 216019 58989
rect 216047 58961 216081 58989
rect 216109 58961 231379 58989
rect 231407 58961 231441 58989
rect 231469 58961 246739 58989
rect 246767 58961 246801 58989
rect 246829 58961 262099 58989
rect 262127 58961 262161 58989
rect 262189 58961 281097 58989
rect 281125 58961 281159 58989
rect 281187 58961 281221 58989
rect 281249 58961 281283 58989
rect 281311 58961 296457 58989
rect 296485 58961 296519 58989
rect 296547 58961 296581 58989
rect 296609 58961 296643 58989
rect 296671 58961 298728 58989
rect 298756 58961 298790 58989
rect 298818 58961 298852 58989
rect 298880 58961 298914 58989
rect 298942 58961 298990 58989
rect -958 58913 298990 58961
rect -958 56175 298990 56223
rect -958 56147 -430 56175
rect -402 56147 -368 56175
rect -340 56147 -306 56175
rect -278 56147 -244 56175
rect -216 56147 2757 56175
rect 2785 56147 2819 56175
rect 2847 56147 2881 56175
rect 2909 56147 2943 56175
rect 2971 56147 18117 56175
rect 18145 56147 18179 56175
rect 18207 56147 18241 56175
rect 18269 56147 18303 56175
rect 18331 56147 33477 56175
rect 33505 56147 33539 56175
rect 33567 56147 33601 56175
rect 33629 56147 33663 56175
rect 33691 56147 48837 56175
rect 48865 56147 48899 56175
rect 48927 56147 48961 56175
rect 48989 56147 49023 56175
rect 49051 56147 64197 56175
rect 64225 56147 64259 56175
rect 64287 56147 64321 56175
rect 64349 56147 64383 56175
rect 64411 56147 79557 56175
rect 79585 56147 79619 56175
rect 79647 56147 79681 56175
rect 79709 56147 79743 56175
rect 79771 56147 94917 56175
rect 94945 56147 94979 56175
rect 95007 56147 95041 56175
rect 95069 56147 95103 56175
rect 95131 56147 110277 56175
rect 110305 56147 110339 56175
rect 110367 56147 110401 56175
rect 110429 56147 110463 56175
rect 110491 56147 125637 56175
rect 125665 56147 125699 56175
rect 125727 56147 125761 56175
rect 125789 56147 125823 56175
rect 125851 56147 140997 56175
rect 141025 56147 141059 56175
rect 141087 56147 141121 56175
rect 141149 56147 141183 56175
rect 141211 56147 156357 56175
rect 156385 56147 156419 56175
rect 156447 56147 156481 56175
rect 156509 56147 156543 56175
rect 156571 56147 162259 56175
rect 162287 56147 162321 56175
rect 162349 56147 177619 56175
rect 177647 56147 177681 56175
rect 177709 56147 192979 56175
rect 193007 56147 193041 56175
rect 193069 56147 208339 56175
rect 208367 56147 208401 56175
rect 208429 56147 223699 56175
rect 223727 56147 223761 56175
rect 223789 56147 239059 56175
rect 239087 56147 239121 56175
rect 239149 56147 254419 56175
rect 254447 56147 254481 56175
rect 254509 56147 269779 56175
rect 269807 56147 269841 56175
rect 269869 56147 279237 56175
rect 279265 56147 279299 56175
rect 279327 56147 279361 56175
rect 279389 56147 279423 56175
rect 279451 56147 294597 56175
rect 294625 56147 294659 56175
rect 294687 56147 294721 56175
rect 294749 56147 294783 56175
rect 294811 56147 298248 56175
rect 298276 56147 298310 56175
rect 298338 56147 298372 56175
rect 298400 56147 298434 56175
rect 298462 56147 298990 56175
rect -958 56113 298990 56147
rect -958 56085 -430 56113
rect -402 56085 -368 56113
rect -340 56085 -306 56113
rect -278 56085 -244 56113
rect -216 56085 2757 56113
rect 2785 56085 2819 56113
rect 2847 56085 2881 56113
rect 2909 56085 2943 56113
rect 2971 56085 18117 56113
rect 18145 56085 18179 56113
rect 18207 56085 18241 56113
rect 18269 56085 18303 56113
rect 18331 56085 33477 56113
rect 33505 56085 33539 56113
rect 33567 56085 33601 56113
rect 33629 56085 33663 56113
rect 33691 56085 48837 56113
rect 48865 56085 48899 56113
rect 48927 56085 48961 56113
rect 48989 56085 49023 56113
rect 49051 56085 64197 56113
rect 64225 56085 64259 56113
rect 64287 56085 64321 56113
rect 64349 56085 64383 56113
rect 64411 56085 79557 56113
rect 79585 56085 79619 56113
rect 79647 56085 79681 56113
rect 79709 56085 79743 56113
rect 79771 56085 94917 56113
rect 94945 56085 94979 56113
rect 95007 56085 95041 56113
rect 95069 56085 95103 56113
rect 95131 56085 110277 56113
rect 110305 56085 110339 56113
rect 110367 56085 110401 56113
rect 110429 56085 110463 56113
rect 110491 56085 125637 56113
rect 125665 56085 125699 56113
rect 125727 56085 125761 56113
rect 125789 56085 125823 56113
rect 125851 56085 140997 56113
rect 141025 56085 141059 56113
rect 141087 56085 141121 56113
rect 141149 56085 141183 56113
rect 141211 56085 156357 56113
rect 156385 56085 156419 56113
rect 156447 56085 156481 56113
rect 156509 56085 156543 56113
rect 156571 56085 162259 56113
rect 162287 56085 162321 56113
rect 162349 56085 177619 56113
rect 177647 56085 177681 56113
rect 177709 56085 192979 56113
rect 193007 56085 193041 56113
rect 193069 56085 208339 56113
rect 208367 56085 208401 56113
rect 208429 56085 223699 56113
rect 223727 56085 223761 56113
rect 223789 56085 239059 56113
rect 239087 56085 239121 56113
rect 239149 56085 254419 56113
rect 254447 56085 254481 56113
rect 254509 56085 269779 56113
rect 269807 56085 269841 56113
rect 269869 56085 279237 56113
rect 279265 56085 279299 56113
rect 279327 56085 279361 56113
rect 279389 56085 279423 56113
rect 279451 56085 294597 56113
rect 294625 56085 294659 56113
rect 294687 56085 294721 56113
rect 294749 56085 294783 56113
rect 294811 56085 298248 56113
rect 298276 56085 298310 56113
rect 298338 56085 298372 56113
rect 298400 56085 298434 56113
rect 298462 56085 298990 56113
rect -958 56051 298990 56085
rect -958 56023 -430 56051
rect -402 56023 -368 56051
rect -340 56023 -306 56051
rect -278 56023 -244 56051
rect -216 56023 2757 56051
rect 2785 56023 2819 56051
rect 2847 56023 2881 56051
rect 2909 56023 2943 56051
rect 2971 56023 18117 56051
rect 18145 56023 18179 56051
rect 18207 56023 18241 56051
rect 18269 56023 18303 56051
rect 18331 56023 33477 56051
rect 33505 56023 33539 56051
rect 33567 56023 33601 56051
rect 33629 56023 33663 56051
rect 33691 56023 48837 56051
rect 48865 56023 48899 56051
rect 48927 56023 48961 56051
rect 48989 56023 49023 56051
rect 49051 56023 64197 56051
rect 64225 56023 64259 56051
rect 64287 56023 64321 56051
rect 64349 56023 64383 56051
rect 64411 56023 79557 56051
rect 79585 56023 79619 56051
rect 79647 56023 79681 56051
rect 79709 56023 79743 56051
rect 79771 56023 94917 56051
rect 94945 56023 94979 56051
rect 95007 56023 95041 56051
rect 95069 56023 95103 56051
rect 95131 56023 110277 56051
rect 110305 56023 110339 56051
rect 110367 56023 110401 56051
rect 110429 56023 110463 56051
rect 110491 56023 125637 56051
rect 125665 56023 125699 56051
rect 125727 56023 125761 56051
rect 125789 56023 125823 56051
rect 125851 56023 140997 56051
rect 141025 56023 141059 56051
rect 141087 56023 141121 56051
rect 141149 56023 141183 56051
rect 141211 56023 156357 56051
rect 156385 56023 156419 56051
rect 156447 56023 156481 56051
rect 156509 56023 156543 56051
rect 156571 56023 162259 56051
rect 162287 56023 162321 56051
rect 162349 56023 177619 56051
rect 177647 56023 177681 56051
rect 177709 56023 192979 56051
rect 193007 56023 193041 56051
rect 193069 56023 208339 56051
rect 208367 56023 208401 56051
rect 208429 56023 223699 56051
rect 223727 56023 223761 56051
rect 223789 56023 239059 56051
rect 239087 56023 239121 56051
rect 239149 56023 254419 56051
rect 254447 56023 254481 56051
rect 254509 56023 269779 56051
rect 269807 56023 269841 56051
rect 269869 56023 279237 56051
rect 279265 56023 279299 56051
rect 279327 56023 279361 56051
rect 279389 56023 279423 56051
rect 279451 56023 294597 56051
rect 294625 56023 294659 56051
rect 294687 56023 294721 56051
rect 294749 56023 294783 56051
rect 294811 56023 298248 56051
rect 298276 56023 298310 56051
rect 298338 56023 298372 56051
rect 298400 56023 298434 56051
rect 298462 56023 298990 56051
rect -958 55989 298990 56023
rect -958 55961 -430 55989
rect -402 55961 -368 55989
rect -340 55961 -306 55989
rect -278 55961 -244 55989
rect -216 55961 2757 55989
rect 2785 55961 2819 55989
rect 2847 55961 2881 55989
rect 2909 55961 2943 55989
rect 2971 55961 18117 55989
rect 18145 55961 18179 55989
rect 18207 55961 18241 55989
rect 18269 55961 18303 55989
rect 18331 55961 33477 55989
rect 33505 55961 33539 55989
rect 33567 55961 33601 55989
rect 33629 55961 33663 55989
rect 33691 55961 48837 55989
rect 48865 55961 48899 55989
rect 48927 55961 48961 55989
rect 48989 55961 49023 55989
rect 49051 55961 64197 55989
rect 64225 55961 64259 55989
rect 64287 55961 64321 55989
rect 64349 55961 64383 55989
rect 64411 55961 79557 55989
rect 79585 55961 79619 55989
rect 79647 55961 79681 55989
rect 79709 55961 79743 55989
rect 79771 55961 94917 55989
rect 94945 55961 94979 55989
rect 95007 55961 95041 55989
rect 95069 55961 95103 55989
rect 95131 55961 110277 55989
rect 110305 55961 110339 55989
rect 110367 55961 110401 55989
rect 110429 55961 110463 55989
rect 110491 55961 125637 55989
rect 125665 55961 125699 55989
rect 125727 55961 125761 55989
rect 125789 55961 125823 55989
rect 125851 55961 140997 55989
rect 141025 55961 141059 55989
rect 141087 55961 141121 55989
rect 141149 55961 141183 55989
rect 141211 55961 156357 55989
rect 156385 55961 156419 55989
rect 156447 55961 156481 55989
rect 156509 55961 156543 55989
rect 156571 55961 162259 55989
rect 162287 55961 162321 55989
rect 162349 55961 177619 55989
rect 177647 55961 177681 55989
rect 177709 55961 192979 55989
rect 193007 55961 193041 55989
rect 193069 55961 208339 55989
rect 208367 55961 208401 55989
rect 208429 55961 223699 55989
rect 223727 55961 223761 55989
rect 223789 55961 239059 55989
rect 239087 55961 239121 55989
rect 239149 55961 254419 55989
rect 254447 55961 254481 55989
rect 254509 55961 269779 55989
rect 269807 55961 269841 55989
rect 269869 55961 279237 55989
rect 279265 55961 279299 55989
rect 279327 55961 279361 55989
rect 279389 55961 279423 55989
rect 279451 55961 294597 55989
rect 294625 55961 294659 55989
rect 294687 55961 294721 55989
rect 294749 55961 294783 55989
rect 294811 55961 298248 55989
rect 298276 55961 298310 55989
rect 298338 55961 298372 55989
rect 298400 55961 298434 55989
rect 298462 55961 298990 55989
rect -958 55913 298990 55961
rect -958 50175 298990 50223
rect -958 50147 -910 50175
rect -882 50147 -848 50175
rect -820 50147 -786 50175
rect -758 50147 -724 50175
rect -696 50147 4617 50175
rect 4645 50147 4679 50175
rect 4707 50147 4741 50175
rect 4769 50147 4803 50175
rect 4831 50147 19977 50175
rect 20005 50147 20039 50175
rect 20067 50147 20101 50175
rect 20129 50147 20163 50175
rect 20191 50147 35337 50175
rect 35365 50147 35399 50175
rect 35427 50147 35461 50175
rect 35489 50147 35523 50175
rect 35551 50147 50697 50175
rect 50725 50147 50759 50175
rect 50787 50147 50821 50175
rect 50849 50147 50883 50175
rect 50911 50147 66057 50175
rect 66085 50147 66119 50175
rect 66147 50147 66181 50175
rect 66209 50147 66243 50175
rect 66271 50147 81417 50175
rect 81445 50147 81479 50175
rect 81507 50147 81541 50175
rect 81569 50147 81603 50175
rect 81631 50147 96777 50175
rect 96805 50147 96839 50175
rect 96867 50147 96901 50175
rect 96929 50147 96963 50175
rect 96991 50147 112137 50175
rect 112165 50147 112199 50175
rect 112227 50147 112261 50175
rect 112289 50147 112323 50175
rect 112351 50147 127497 50175
rect 127525 50147 127559 50175
rect 127587 50147 127621 50175
rect 127649 50147 127683 50175
rect 127711 50147 142857 50175
rect 142885 50147 142919 50175
rect 142947 50147 142981 50175
rect 143009 50147 143043 50175
rect 143071 50147 158217 50175
rect 158245 50147 158279 50175
rect 158307 50147 158341 50175
rect 158369 50147 158403 50175
rect 158431 50147 169939 50175
rect 169967 50147 170001 50175
rect 170029 50147 185299 50175
rect 185327 50147 185361 50175
rect 185389 50147 200659 50175
rect 200687 50147 200721 50175
rect 200749 50147 216019 50175
rect 216047 50147 216081 50175
rect 216109 50147 231379 50175
rect 231407 50147 231441 50175
rect 231469 50147 246739 50175
rect 246767 50147 246801 50175
rect 246829 50147 262099 50175
rect 262127 50147 262161 50175
rect 262189 50147 281097 50175
rect 281125 50147 281159 50175
rect 281187 50147 281221 50175
rect 281249 50147 281283 50175
rect 281311 50147 296457 50175
rect 296485 50147 296519 50175
rect 296547 50147 296581 50175
rect 296609 50147 296643 50175
rect 296671 50147 298728 50175
rect 298756 50147 298790 50175
rect 298818 50147 298852 50175
rect 298880 50147 298914 50175
rect 298942 50147 298990 50175
rect -958 50113 298990 50147
rect -958 50085 -910 50113
rect -882 50085 -848 50113
rect -820 50085 -786 50113
rect -758 50085 -724 50113
rect -696 50085 4617 50113
rect 4645 50085 4679 50113
rect 4707 50085 4741 50113
rect 4769 50085 4803 50113
rect 4831 50085 19977 50113
rect 20005 50085 20039 50113
rect 20067 50085 20101 50113
rect 20129 50085 20163 50113
rect 20191 50085 35337 50113
rect 35365 50085 35399 50113
rect 35427 50085 35461 50113
rect 35489 50085 35523 50113
rect 35551 50085 50697 50113
rect 50725 50085 50759 50113
rect 50787 50085 50821 50113
rect 50849 50085 50883 50113
rect 50911 50085 66057 50113
rect 66085 50085 66119 50113
rect 66147 50085 66181 50113
rect 66209 50085 66243 50113
rect 66271 50085 81417 50113
rect 81445 50085 81479 50113
rect 81507 50085 81541 50113
rect 81569 50085 81603 50113
rect 81631 50085 96777 50113
rect 96805 50085 96839 50113
rect 96867 50085 96901 50113
rect 96929 50085 96963 50113
rect 96991 50085 112137 50113
rect 112165 50085 112199 50113
rect 112227 50085 112261 50113
rect 112289 50085 112323 50113
rect 112351 50085 127497 50113
rect 127525 50085 127559 50113
rect 127587 50085 127621 50113
rect 127649 50085 127683 50113
rect 127711 50085 142857 50113
rect 142885 50085 142919 50113
rect 142947 50085 142981 50113
rect 143009 50085 143043 50113
rect 143071 50085 158217 50113
rect 158245 50085 158279 50113
rect 158307 50085 158341 50113
rect 158369 50085 158403 50113
rect 158431 50085 169939 50113
rect 169967 50085 170001 50113
rect 170029 50085 185299 50113
rect 185327 50085 185361 50113
rect 185389 50085 200659 50113
rect 200687 50085 200721 50113
rect 200749 50085 216019 50113
rect 216047 50085 216081 50113
rect 216109 50085 231379 50113
rect 231407 50085 231441 50113
rect 231469 50085 246739 50113
rect 246767 50085 246801 50113
rect 246829 50085 262099 50113
rect 262127 50085 262161 50113
rect 262189 50085 281097 50113
rect 281125 50085 281159 50113
rect 281187 50085 281221 50113
rect 281249 50085 281283 50113
rect 281311 50085 296457 50113
rect 296485 50085 296519 50113
rect 296547 50085 296581 50113
rect 296609 50085 296643 50113
rect 296671 50085 298728 50113
rect 298756 50085 298790 50113
rect 298818 50085 298852 50113
rect 298880 50085 298914 50113
rect 298942 50085 298990 50113
rect -958 50051 298990 50085
rect -958 50023 -910 50051
rect -882 50023 -848 50051
rect -820 50023 -786 50051
rect -758 50023 -724 50051
rect -696 50023 4617 50051
rect 4645 50023 4679 50051
rect 4707 50023 4741 50051
rect 4769 50023 4803 50051
rect 4831 50023 19977 50051
rect 20005 50023 20039 50051
rect 20067 50023 20101 50051
rect 20129 50023 20163 50051
rect 20191 50023 35337 50051
rect 35365 50023 35399 50051
rect 35427 50023 35461 50051
rect 35489 50023 35523 50051
rect 35551 50023 50697 50051
rect 50725 50023 50759 50051
rect 50787 50023 50821 50051
rect 50849 50023 50883 50051
rect 50911 50023 66057 50051
rect 66085 50023 66119 50051
rect 66147 50023 66181 50051
rect 66209 50023 66243 50051
rect 66271 50023 81417 50051
rect 81445 50023 81479 50051
rect 81507 50023 81541 50051
rect 81569 50023 81603 50051
rect 81631 50023 96777 50051
rect 96805 50023 96839 50051
rect 96867 50023 96901 50051
rect 96929 50023 96963 50051
rect 96991 50023 112137 50051
rect 112165 50023 112199 50051
rect 112227 50023 112261 50051
rect 112289 50023 112323 50051
rect 112351 50023 127497 50051
rect 127525 50023 127559 50051
rect 127587 50023 127621 50051
rect 127649 50023 127683 50051
rect 127711 50023 142857 50051
rect 142885 50023 142919 50051
rect 142947 50023 142981 50051
rect 143009 50023 143043 50051
rect 143071 50023 158217 50051
rect 158245 50023 158279 50051
rect 158307 50023 158341 50051
rect 158369 50023 158403 50051
rect 158431 50023 169939 50051
rect 169967 50023 170001 50051
rect 170029 50023 185299 50051
rect 185327 50023 185361 50051
rect 185389 50023 200659 50051
rect 200687 50023 200721 50051
rect 200749 50023 216019 50051
rect 216047 50023 216081 50051
rect 216109 50023 231379 50051
rect 231407 50023 231441 50051
rect 231469 50023 246739 50051
rect 246767 50023 246801 50051
rect 246829 50023 262099 50051
rect 262127 50023 262161 50051
rect 262189 50023 281097 50051
rect 281125 50023 281159 50051
rect 281187 50023 281221 50051
rect 281249 50023 281283 50051
rect 281311 50023 296457 50051
rect 296485 50023 296519 50051
rect 296547 50023 296581 50051
rect 296609 50023 296643 50051
rect 296671 50023 298728 50051
rect 298756 50023 298790 50051
rect 298818 50023 298852 50051
rect 298880 50023 298914 50051
rect 298942 50023 298990 50051
rect -958 49989 298990 50023
rect -958 49961 -910 49989
rect -882 49961 -848 49989
rect -820 49961 -786 49989
rect -758 49961 -724 49989
rect -696 49961 4617 49989
rect 4645 49961 4679 49989
rect 4707 49961 4741 49989
rect 4769 49961 4803 49989
rect 4831 49961 19977 49989
rect 20005 49961 20039 49989
rect 20067 49961 20101 49989
rect 20129 49961 20163 49989
rect 20191 49961 35337 49989
rect 35365 49961 35399 49989
rect 35427 49961 35461 49989
rect 35489 49961 35523 49989
rect 35551 49961 50697 49989
rect 50725 49961 50759 49989
rect 50787 49961 50821 49989
rect 50849 49961 50883 49989
rect 50911 49961 66057 49989
rect 66085 49961 66119 49989
rect 66147 49961 66181 49989
rect 66209 49961 66243 49989
rect 66271 49961 81417 49989
rect 81445 49961 81479 49989
rect 81507 49961 81541 49989
rect 81569 49961 81603 49989
rect 81631 49961 96777 49989
rect 96805 49961 96839 49989
rect 96867 49961 96901 49989
rect 96929 49961 96963 49989
rect 96991 49961 112137 49989
rect 112165 49961 112199 49989
rect 112227 49961 112261 49989
rect 112289 49961 112323 49989
rect 112351 49961 127497 49989
rect 127525 49961 127559 49989
rect 127587 49961 127621 49989
rect 127649 49961 127683 49989
rect 127711 49961 142857 49989
rect 142885 49961 142919 49989
rect 142947 49961 142981 49989
rect 143009 49961 143043 49989
rect 143071 49961 158217 49989
rect 158245 49961 158279 49989
rect 158307 49961 158341 49989
rect 158369 49961 158403 49989
rect 158431 49961 169939 49989
rect 169967 49961 170001 49989
rect 170029 49961 185299 49989
rect 185327 49961 185361 49989
rect 185389 49961 200659 49989
rect 200687 49961 200721 49989
rect 200749 49961 216019 49989
rect 216047 49961 216081 49989
rect 216109 49961 231379 49989
rect 231407 49961 231441 49989
rect 231469 49961 246739 49989
rect 246767 49961 246801 49989
rect 246829 49961 262099 49989
rect 262127 49961 262161 49989
rect 262189 49961 281097 49989
rect 281125 49961 281159 49989
rect 281187 49961 281221 49989
rect 281249 49961 281283 49989
rect 281311 49961 296457 49989
rect 296485 49961 296519 49989
rect 296547 49961 296581 49989
rect 296609 49961 296643 49989
rect 296671 49961 298728 49989
rect 298756 49961 298790 49989
rect 298818 49961 298852 49989
rect 298880 49961 298914 49989
rect 298942 49961 298990 49989
rect -958 49913 298990 49961
rect -958 47175 298990 47223
rect -958 47147 -430 47175
rect -402 47147 -368 47175
rect -340 47147 -306 47175
rect -278 47147 -244 47175
rect -216 47147 2757 47175
rect 2785 47147 2819 47175
rect 2847 47147 2881 47175
rect 2909 47147 2943 47175
rect 2971 47147 18117 47175
rect 18145 47147 18179 47175
rect 18207 47147 18241 47175
rect 18269 47147 18303 47175
rect 18331 47147 33477 47175
rect 33505 47147 33539 47175
rect 33567 47147 33601 47175
rect 33629 47147 33663 47175
rect 33691 47147 48837 47175
rect 48865 47147 48899 47175
rect 48927 47147 48961 47175
rect 48989 47147 49023 47175
rect 49051 47147 64197 47175
rect 64225 47147 64259 47175
rect 64287 47147 64321 47175
rect 64349 47147 64383 47175
rect 64411 47147 79557 47175
rect 79585 47147 79619 47175
rect 79647 47147 79681 47175
rect 79709 47147 79743 47175
rect 79771 47147 94917 47175
rect 94945 47147 94979 47175
rect 95007 47147 95041 47175
rect 95069 47147 95103 47175
rect 95131 47147 110277 47175
rect 110305 47147 110339 47175
rect 110367 47147 110401 47175
rect 110429 47147 110463 47175
rect 110491 47147 125637 47175
rect 125665 47147 125699 47175
rect 125727 47147 125761 47175
rect 125789 47147 125823 47175
rect 125851 47147 140997 47175
rect 141025 47147 141059 47175
rect 141087 47147 141121 47175
rect 141149 47147 141183 47175
rect 141211 47147 156357 47175
rect 156385 47147 156419 47175
rect 156447 47147 156481 47175
rect 156509 47147 156543 47175
rect 156571 47147 162259 47175
rect 162287 47147 162321 47175
rect 162349 47147 177619 47175
rect 177647 47147 177681 47175
rect 177709 47147 192979 47175
rect 193007 47147 193041 47175
rect 193069 47147 208339 47175
rect 208367 47147 208401 47175
rect 208429 47147 223699 47175
rect 223727 47147 223761 47175
rect 223789 47147 239059 47175
rect 239087 47147 239121 47175
rect 239149 47147 254419 47175
rect 254447 47147 254481 47175
rect 254509 47147 269779 47175
rect 269807 47147 269841 47175
rect 269869 47147 279237 47175
rect 279265 47147 279299 47175
rect 279327 47147 279361 47175
rect 279389 47147 279423 47175
rect 279451 47147 294597 47175
rect 294625 47147 294659 47175
rect 294687 47147 294721 47175
rect 294749 47147 294783 47175
rect 294811 47147 298248 47175
rect 298276 47147 298310 47175
rect 298338 47147 298372 47175
rect 298400 47147 298434 47175
rect 298462 47147 298990 47175
rect -958 47113 298990 47147
rect -958 47085 -430 47113
rect -402 47085 -368 47113
rect -340 47085 -306 47113
rect -278 47085 -244 47113
rect -216 47085 2757 47113
rect 2785 47085 2819 47113
rect 2847 47085 2881 47113
rect 2909 47085 2943 47113
rect 2971 47085 18117 47113
rect 18145 47085 18179 47113
rect 18207 47085 18241 47113
rect 18269 47085 18303 47113
rect 18331 47085 33477 47113
rect 33505 47085 33539 47113
rect 33567 47085 33601 47113
rect 33629 47085 33663 47113
rect 33691 47085 48837 47113
rect 48865 47085 48899 47113
rect 48927 47085 48961 47113
rect 48989 47085 49023 47113
rect 49051 47085 64197 47113
rect 64225 47085 64259 47113
rect 64287 47085 64321 47113
rect 64349 47085 64383 47113
rect 64411 47085 79557 47113
rect 79585 47085 79619 47113
rect 79647 47085 79681 47113
rect 79709 47085 79743 47113
rect 79771 47085 94917 47113
rect 94945 47085 94979 47113
rect 95007 47085 95041 47113
rect 95069 47085 95103 47113
rect 95131 47085 110277 47113
rect 110305 47085 110339 47113
rect 110367 47085 110401 47113
rect 110429 47085 110463 47113
rect 110491 47085 125637 47113
rect 125665 47085 125699 47113
rect 125727 47085 125761 47113
rect 125789 47085 125823 47113
rect 125851 47085 140997 47113
rect 141025 47085 141059 47113
rect 141087 47085 141121 47113
rect 141149 47085 141183 47113
rect 141211 47085 156357 47113
rect 156385 47085 156419 47113
rect 156447 47085 156481 47113
rect 156509 47085 156543 47113
rect 156571 47085 162259 47113
rect 162287 47085 162321 47113
rect 162349 47085 177619 47113
rect 177647 47085 177681 47113
rect 177709 47085 192979 47113
rect 193007 47085 193041 47113
rect 193069 47085 208339 47113
rect 208367 47085 208401 47113
rect 208429 47085 223699 47113
rect 223727 47085 223761 47113
rect 223789 47085 239059 47113
rect 239087 47085 239121 47113
rect 239149 47085 254419 47113
rect 254447 47085 254481 47113
rect 254509 47085 269779 47113
rect 269807 47085 269841 47113
rect 269869 47085 279237 47113
rect 279265 47085 279299 47113
rect 279327 47085 279361 47113
rect 279389 47085 279423 47113
rect 279451 47085 294597 47113
rect 294625 47085 294659 47113
rect 294687 47085 294721 47113
rect 294749 47085 294783 47113
rect 294811 47085 298248 47113
rect 298276 47085 298310 47113
rect 298338 47085 298372 47113
rect 298400 47085 298434 47113
rect 298462 47085 298990 47113
rect -958 47051 298990 47085
rect -958 47023 -430 47051
rect -402 47023 -368 47051
rect -340 47023 -306 47051
rect -278 47023 -244 47051
rect -216 47023 2757 47051
rect 2785 47023 2819 47051
rect 2847 47023 2881 47051
rect 2909 47023 2943 47051
rect 2971 47023 18117 47051
rect 18145 47023 18179 47051
rect 18207 47023 18241 47051
rect 18269 47023 18303 47051
rect 18331 47023 33477 47051
rect 33505 47023 33539 47051
rect 33567 47023 33601 47051
rect 33629 47023 33663 47051
rect 33691 47023 48837 47051
rect 48865 47023 48899 47051
rect 48927 47023 48961 47051
rect 48989 47023 49023 47051
rect 49051 47023 64197 47051
rect 64225 47023 64259 47051
rect 64287 47023 64321 47051
rect 64349 47023 64383 47051
rect 64411 47023 79557 47051
rect 79585 47023 79619 47051
rect 79647 47023 79681 47051
rect 79709 47023 79743 47051
rect 79771 47023 94917 47051
rect 94945 47023 94979 47051
rect 95007 47023 95041 47051
rect 95069 47023 95103 47051
rect 95131 47023 110277 47051
rect 110305 47023 110339 47051
rect 110367 47023 110401 47051
rect 110429 47023 110463 47051
rect 110491 47023 125637 47051
rect 125665 47023 125699 47051
rect 125727 47023 125761 47051
rect 125789 47023 125823 47051
rect 125851 47023 140997 47051
rect 141025 47023 141059 47051
rect 141087 47023 141121 47051
rect 141149 47023 141183 47051
rect 141211 47023 156357 47051
rect 156385 47023 156419 47051
rect 156447 47023 156481 47051
rect 156509 47023 156543 47051
rect 156571 47023 162259 47051
rect 162287 47023 162321 47051
rect 162349 47023 177619 47051
rect 177647 47023 177681 47051
rect 177709 47023 192979 47051
rect 193007 47023 193041 47051
rect 193069 47023 208339 47051
rect 208367 47023 208401 47051
rect 208429 47023 223699 47051
rect 223727 47023 223761 47051
rect 223789 47023 239059 47051
rect 239087 47023 239121 47051
rect 239149 47023 254419 47051
rect 254447 47023 254481 47051
rect 254509 47023 269779 47051
rect 269807 47023 269841 47051
rect 269869 47023 279237 47051
rect 279265 47023 279299 47051
rect 279327 47023 279361 47051
rect 279389 47023 279423 47051
rect 279451 47023 294597 47051
rect 294625 47023 294659 47051
rect 294687 47023 294721 47051
rect 294749 47023 294783 47051
rect 294811 47023 298248 47051
rect 298276 47023 298310 47051
rect 298338 47023 298372 47051
rect 298400 47023 298434 47051
rect 298462 47023 298990 47051
rect -958 46989 298990 47023
rect -958 46961 -430 46989
rect -402 46961 -368 46989
rect -340 46961 -306 46989
rect -278 46961 -244 46989
rect -216 46961 2757 46989
rect 2785 46961 2819 46989
rect 2847 46961 2881 46989
rect 2909 46961 2943 46989
rect 2971 46961 18117 46989
rect 18145 46961 18179 46989
rect 18207 46961 18241 46989
rect 18269 46961 18303 46989
rect 18331 46961 33477 46989
rect 33505 46961 33539 46989
rect 33567 46961 33601 46989
rect 33629 46961 33663 46989
rect 33691 46961 48837 46989
rect 48865 46961 48899 46989
rect 48927 46961 48961 46989
rect 48989 46961 49023 46989
rect 49051 46961 64197 46989
rect 64225 46961 64259 46989
rect 64287 46961 64321 46989
rect 64349 46961 64383 46989
rect 64411 46961 79557 46989
rect 79585 46961 79619 46989
rect 79647 46961 79681 46989
rect 79709 46961 79743 46989
rect 79771 46961 94917 46989
rect 94945 46961 94979 46989
rect 95007 46961 95041 46989
rect 95069 46961 95103 46989
rect 95131 46961 110277 46989
rect 110305 46961 110339 46989
rect 110367 46961 110401 46989
rect 110429 46961 110463 46989
rect 110491 46961 125637 46989
rect 125665 46961 125699 46989
rect 125727 46961 125761 46989
rect 125789 46961 125823 46989
rect 125851 46961 140997 46989
rect 141025 46961 141059 46989
rect 141087 46961 141121 46989
rect 141149 46961 141183 46989
rect 141211 46961 156357 46989
rect 156385 46961 156419 46989
rect 156447 46961 156481 46989
rect 156509 46961 156543 46989
rect 156571 46961 162259 46989
rect 162287 46961 162321 46989
rect 162349 46961 177619 46989
rect 177647 46961 177681 46989
rect 177709 46961 192979 46989
rect 193007 46961 193041 46989
rect 193069 46961 208339 46989
rect 208367 46961 208401 46989
rect 208429 46961 223699 46989
rect 223727 46961 223761 46989
rect 223789 46961 239059 46989
rect 239087 46961 239121 46989
rect 239149 46961 254419 46989
rect 254447 46961 254481 46989
rect 254509 46961 269779 46989
rect 269807 46961 269841 46989
rect 269869 46961 279237 46989
rect 279265 46961 279299 46989
rect 279327 46961 279361 46989
rect 279389 46961 279423 46989
rect 279451 46961 294597 46989
rect 294625 46961 294659 46989
rect 294687 46961 294721 46989
rect 294749 46961 294783 46989
rect 294811 46961 298248 46989
rect 298276 46961 298310 46989
rect 298338 46961 298372 46989
rect 298400 46961 298434 46989
rect 298462 46961 298990 46989
rect -958 46913 298990 46961
rect -958 41175 298990 41223
rect -958 41147 -910 41175
rect -882 41147 -848 41175
rect -820 41147 -786 41175
rect -758 41147 -724 41175
rect -696 41147 4617 41175
rect 4645 41147 4679 41175
rect 4707 41147 4741 41175
rect 4769 41147 4803 41175
rect 4831 41147 19977 41175
rect 20005 41147 20039 41175
rect 20067 41147 20101 41175
rect 20129 41147 20163 41175
rect 20191 41147 35337 41175
rect 35365 41147 35399 41175
rect 35427 41147 35461 41175
rect 35489 41147 35523 41175
rect 35551 41147 50697 41175
rect 50725 41147 50759 41175
rect 50787 41147 50821 41175
rect 50849 41147 50883 41175
rect 50911 41147 66057 41175
rect 66085 41147 66119 41175
rect 66147 41147 66181 41175
rect 66209 41147 66243 41175
rect 66271 41147 81417 41175
rect 81445 41147 81479 41175
rect 81507 41147 81541 41175
rect 81569 41147 81603 41175
rect 81631 41147 96777 41175
rect 96805 41147 96839 41175
rect 96867 41147 96901 41175
rect 96929 41147 96963 41175
rect 96991 41147 112137 41175
rect 112165 41147 112199 41175
rect 112227 41147 112261 41175
rect 112289 41147 112323 41175
rect 112351 41147 127497 41175
rect 127525 41147 127559 41175
rect 127587 41147 127621 41175
rect 127649 41147 127683 41175
rect 127711 41147 142857 41175
rect 142885 41147 142919 41175
rect 142947 41147 142981 41175
rect 143009 41147 143043 41175
rect 143071 41147 158217 41175
rect 158245 41147 158279 41175
rect 158307 41147 158341 41175
rect 158369 41147 158403 41175
rect 158431 41147 169939 41175
rect 169967 41147 170001 41175
rect 170029 41147 185299 41175
rect 185327 41147 185361 41175
rect 185389 41147 200659 41175
rect 200687 41147 200721 41175
rect 200749 41147 216019 41175
rect 216047 41147 216081 41175
rect 216109 41147 231379 41175
rect 231407 41147 231441 41175
rect 231469 41147 246739 41175
rect 246767 41147 246801 41175
rect 246829 41147 262099 41175
rect 262127 41147 262161 41175
rect 262189 41147 281097 41175
rect 281125 41147 281159 41175
rect 281187 41147 281221 41175
rect 281249 41147 281283 41175
rect 281311 41147 296457 41175
rect 296485 41147 296519 41175
rect 296547 41147 296581 41175
rect 296609 41147 296643 41175
rect 296671 41147 298728 41175
rect 298756 41147 298790 41175
rect 298818 41147 298852 41175
rect 298880 41147 298914 41175
rect 298942 41147 298990 41175
rect -958 41113 298990 41147
rect -958 41085 -910 41113
rect -882 41085 -848 41113
rect -820 41085 -786 41113
rect -758 41085 -724 41113
rect -696 41085 4617 41113
rect 4645 41085 4679 41113
rect 4707 41085 4741 41113
rect 4769 41085 4803 41113
rect 4831 41085 19977 41113
rect 20005 41085 20039 41113
rect 20067 41085 20101 41113
rect 20129 41085 20163 41113
rect 20191 41085 35337 41113
rect 35365 41085 35399 41113
rect 35427 41085 35461 41113
rect 35489 41085 35523 41113
rect 35551 41085 50697 41113
rect 50725 41085 50759 41113
rect 50787 41085 50821 41113
rect 50849 41085 50883 41113
rect 50911 41085 66057 41113
rect 66085 41085 66119 41113
rect 66147 41085 66181 41113
rect 66209 41085 66243 41113
rect 66271 41085 81417 41113
rect 81445 41085 81479 41113
rect 81507 41085 81541 41113
rect 81569 41085 81603 41113
rect 81631 41085 96777 41113
rect 96805 41085 96839 41113
rect 96867 41085 96901 41113
rect 96929 41085 96963 41113
rect 96991 41085 112137 41113
rect 112165 41085 112199 41113
rect 112227 41085 112261 41113
rect 112289 41085 112323 41113
rect 112351 41085 127497 41113
rect 127525 41085 127559 41113
rect 127587 41085 127621 41113
rect 127649 41085 127683 41113
rect 127711 41085 142857 41113
rect 142885 41085 142919 41113
rect 142947 41085 142981 41113
rect 143009 41085 143043 41113
rect 143071 41085 158217 41113
rect 158245 41085 158279 41113
rect 158307 41085 158341 41113
rect 158369 41085 158403 41113
rect 158431 41085 169939 41113
rect 169967 41085 170001 41113
rect 170029 41085 185299 41113
rect 185327 41085 185361 41113
rect 185389 41085 200659 41113
rect 200687 41085 200721 41113
rect 200749 41085 216019 41113
rect 216047 41085 216081 41113
rect 216109 41085 231379 41113
rect 231407 41085 231441 41113
rect 231469 41085 246739 41113
rect 246767 41085 246801 41113
rect 246829 41085 262099 41113
rect 262127 41085 262161 41113
rect 262189 41085 281097 41113
rect 281125 41085 281159 41113
rect 281187 41085 281221 41113
rect 281249 41085 281283 41113
rect 281311 41085 296457 41113
rect 296485 41085 296519 41113
rect 296547 41085 296581 41113
rect 296609 41085 296643 41113
rect 296671 41085 298728 41113
rect 298756 41085 298790 41113
rect 298818 41085 298852 41113
rect 298880 41085 298914 41113
rect 298942 41085 298990 41113
rect -958 41051 298990 41085
rect -958 41023 -910 41051
rect -882 41023 -848 41051
rect -820 41023 -786 41051
rect -758 41023 -724 41051
rect -696 41023 4617 41051
rect 4645 41023 4679 41051
rect 4707 41023 4741 41051
rect 4769 41023 4803 41051
rect 4831 41023 19977 41051
rect 20005 41023 20039 41051
rect 20067 41023 20101 41051
rect 20129 41023 20163 41051
rect 20191 41023 35337 41051
rect 35365 41023 35399 41051
rect 35427 41023 35461 41051
rect 35489 41023 35523 41051
rect 35551 41023 50697 41051
rect 50725 41023 50759 41051
rect 50787 41023 50821 41051
rect 50849 41023 50883 41051
rect 50911 41023 66057 41051
rect 66085 41023 66119 41051
rect 66147 41023 66181 41051
rect 66209 41023 66243 41051
rect 66271 41023 81417 41051
rect 81445 41023 81479 41051
rect 81507 41023 81541 41051
rect 81569 41023 81603 41051
rect 81631 41023 96777 41051
rect 96805 41023 96839 41051
rect 96867 41023 96901 41051
rect 96929 41023 96963 41051
rect 96991 41023 112137 41051
rect 112165 41023 112199 41051
rect 112227 41023 112261 41051
rect 112289 41023 112323 41051
rect 112351 41023 127497 41051
rect 127525 41023 127559 41051
rect 127587 41023 127621 41051
rect 127649 41023 127683 41051
rect 127711 41023 142857 41051
rect 142885 41023 142919 41051
rect 142947 41023 142981 41051
rect 143009 41023 143043 41051
rect 143071 41023 158217 41051
rect 158245 41023 158279 41051
rect 158307 41023 158341 41051
rect 158369 41023 158403 41051
rect 158431 41023 169939 41051
rect 169967 41023 170001 41051
rect 170029 41023 185299 41051
rect 185327 41023 185361 41051
rect 185389 41023 200659 41051
rect 200687 41023 200721 41051
rect 200749 41023 216019 41051
rect 216047 41023 216081 41051
rect 216109 41023 231379 41051
rect 231407 41023 231441 41051
rect 231469 41023 246739 41051
rect 246767 41023 246801 41051
rect 246829 41023 262099 41051
rect 262127 41023 262161 41051
rect 262189 41023 281097 41051
rect 281125 41023 281159 41051
rect 281187 41023 281221 41051
rect 281249 41023 281283 41051
rect 281311 41023 296457 41051
rect 296485 41023 296519 41051
rect 296547 41023 296581 41051
rect 296609 41023 296643 41051
rect 296671 41023 298728 41051
rect 298756 41023 298790 41051
rect 298818 41023 298852 41051
rect 298880 41023 298914 41051
rect 298942 41023 298990 41051
rect -958 40989 298990 41023
rect -958 40961 -910 40989
rect -882 40961 -848 40989
rect -820 40961 -786 40989
rect -758 40961 -724 40989
rect -696 40961 4617 40989
rect 4645 40961 4679 40989
rect 4707 40961 4741 40989
rect 4769 40961 4803 40989
rect 4831 40961 19977 40989
rect 20005 40961 20039 40989
rect 20067 40961 20101 40989
rect 20129 40961 20163 40989
rect 20191 40961 35337 40989
rect 35365 40961 35399 40989
rect 35427 40961 35461 40989
rect 35489 40961 35523 40989
rect 35551 40961 50697 40989
rect 50725 40961 50759 40989
rect 50787 40961 50821 40989
rect 50849 40961 50883 40989
rect 50911 40961 66057 40989
rect 66085 40961 66119 40989
rect 66147 40961 66181 40989
rect 66209 40961 66243 40989
rect 66271 40961 81417 40989
rect 81445 40961 81479 40989
rect 81507 40961 81541 40989
rect 81569 40961 81603 40989
rect 81631 40961 96777 40989
rect 96805 40961 96839 40989
rect 96867 40961 96901 40989
rect 96929 40961 96963 40989
rect 96991 40961 112137 40989
rect 112165 40961 112199 40989
rect 112227 40961 112261 40989
rect 112289 40961 112323 40989
rect 112351 40961 127497 40989
rect 127525 40961 127559 40989
rect 127587 40961 127621 40989
rect 127649 40961 127683 40989
rect 127711 40961 142857 40989
rect 142885 40961 142919 40989
rect 142947 40961 142981 40989
rect 143009 40961 143043 40989
rect 143071 40961 158217 40989
rect 158245 40961 158279 40989
rect 158307 40961 158341 40989
rect 158369 40961 158403 40989
rect 158431 40961 169939 40989
rect 169967 40961 170001 40989
rect 170029 40961 185299 40989
rect 185327 40961 185361 40989
rect 185389 40961 200659 40989
rect 200687 40961 200721 40989
rect 200749 40961 216019 40989
rect 216047 40961 216081 40989
rect 216109 40961 231379 40989
rect 231407 40961 231441 40989
rect 231469 40961 246739 40989
rect 246767 40961 246801 40989
rect 246829 40961 262099 40989
rect 262127 40961 262161 40989
rect 262189 40961 281097 40989
rect 281125 40961 281159 40989
rect 281187 40961 281221 40989
rect 281249 40961 281283 40989
rect 281311 40961 296457 40989
rect 296485 40961 296519 40989
rect 296547 40961 296581 40989
rect 296609 40961 296643 40989
rect 296671 40961 298728 40989
rect 298756 40961 298790 40989
rect 298818 40961 298852 40989
rect 298880 40961 298914 40989
rect 298942 40961 298990 40989
rect -958 40913 298990 40961
rect -958 38175 298990 38223
rect -958 38147 -430 38175
rect -402 38147 -368 38175
rect -340 38147 -306 38175
rect -278 38147 -244 38175
rect -216 38147 2757 38175
rect 2785 38147 2819 38175
rect 2847 38147 2881 38175
rect 2909 38147 2943 38175
rect 2971 38147 18117 38175
rect 18145 38147 18179 38175
rect 18207 38147 18241 38175
rect 18269 38147 18303 38175
rect 18331 38147 33477 38175
rect 33505 38147 33539 38175
rect 33567 38147 33601 38175
rect 33629 38147 33663 38175
rect 33691 38147 48837 38175
rect 48865 38147 48899 38175
rect 48927 38147 48961 38175
rect 48989 38147 49023 38175
rect 49051 38147 64197 38175
rect 64225 38147 64259 38175
rect 64287 38147 64321 38175
rect 64349 38147 64383 38175
rect 64411 38147 79557 38175
rect 79585 38147 79619 38175
rect 79647 38147 79681 38175
rect 79709 38147 79743 38175
rect 79771 38147 94917 38175
rect 94945 38147 94979 38175
rect 95007 38147 95041 38175
rect 95069 38147 95103 38175
rect 95131 38147 110277 38175
rect 110305 38147 110339 38175
rect 110367 38147 110401 38175
rect 110429 38147 110463 38175
rect 110491 38147 125637 38175
rect 125665 38147 125699 38175
rect 125727 38147 125761 38175
rect 125789 38147 125823 38175
rect 125851 38147 140997 38175
rect 141025 38147 141059 38175
rect 141087 38147 141121 38175
rect 141149 38147 141183 38175
rect 141211 38147 156357 38175
rect 156385 38147 156419 38175
rect 156447 38147 156481 38175
rect 156509 38147 156543 38175
rect 156571 38147 162259 38175
rect 162287 38147 162321 38175
rect 162349 38147 177619 38175
rect 177647 38147 177681 38175
rect 177709 38147 192979 38175
rect 193007 38147 193041 38175
rect 193069 38147 208339 38175
rect 208367 38147 208401 38175
rect 208429 38147 223699 38175
rect 223727 38147 223761 38175
rect 223789 38147 239059 38175
rect 239087 38147 239121 38175
rect 239149 38147 254419 38175
rect 254447 38147 254481 38175
rect 254509 38147 269779 38175
rect 269807 38147 269841 38175
rect 269869 38147 279237 38175
rect 279265 38147 279299 38175
rect 279327 38147 279361 38175
rect 279389 38147 279423 38175
rect 279451 38147 294597 38175
rect 294625 38147 294659 38175
rect 294687 38147 294721 38175
rect 294749 38147 294783 38175
rect 294811 38147 298248 38175
rect 298276 38147 298310 38175
rect 298338 38147 298372 38175
rect 298400 38147 298434 38175
rect 298462 38147 298990 38175
rect -958 38113 298990 38147
rect -958 38085 -430 38113
rect -402 38085 -368 38113
rect -340 38085 -306 38113
rect -278 38085 -244 38113
rect -216 38085 2757 38113
rect 2785 38085 2819 38113
rect 2847 38085 2881 38113
rect 2909 38085 2943 38113
rect 2971 38085 18117 38113
rect 18145 38085 18179 38113
rect 18207 38085 18241 38113
rect 18269 38085 18303 38113
rect 18331 38085 33477 38113
rect 33505 38085 33539 38113
rect 33567 38085 33601 38113
rect 33629 38085 33663 38113
rect 33691 38085 48837 38113
rect 48865 38085 48899 38113
rect 48927 38085 48961 38113
rect 48989 38085 49023 38113
rect 49051 38085 64197 38113
rect 64225 38085 64259 38113
rect 64287 38085 64321 38113
rect 64349 38085 64383 38113
rect 64411 38085 79557 38113
rect 79585 38085 79619 38113
rect 79647 38085 79681 38113
rect 79709 38085 79743 38113
rect 79771 38085 94917 38113
rect 94945 38085 94979 38113
rect 95007 38085 95041 38113
rect 95069 38085 95103 38113
rect 95131 38085 110277 38113
rect 110305 38085 110339 38113
rect 110367 38085 110401 38113
rect 110429 38085 110463 38113
rect 110491 38085 125637 38113
rect 125665 38085 125699 38113
rect 125727 38085 125761 38113
rect 125789 38085 125823 38113
rect 125851 38085 140997 38113
rect 141025 38085 141059 38113
rect 141087 38085 141121 38113
rect 141149 38085 141183 38113
rect 141211 38085 156357 38113
rect 156385 38085 156419 38113
rect 156447 38085 156481 38113
rect 156509 38085 156543 38113
rect 156571 38085 162259 38113
rect 162287 38085 162321 38113
rect 162349 38085 177619 38113
rect 177647 38085 177681 38113
rect 177709 38085 192979 38113
rect 193007 38085 193041 38113
rect 193069 38085 208339 38113
rect 208367 38085 208401 38113
rect 208429 38085 223699 38113
rect 223727 38085 223761 38113
rect 223789 38085 239059 38113
rect 239087 38085 239121 38113
rect 239149 38085 254419 38113
rect 254447 38085 254481 38113
rect 254509 38085 269779 38113
rect 269807 38085 269841 38113
rect 269869 38085 279237 38113
rect 279265 38085 279299 38113
rect 279327 38085 279361 38113
rect 279389 38085 279423 38113
rect 279451 38085 294597 38113
rect 294625 38085 294659 38113
rect 294687 38085 294721 38113
rect 294749 38085 294783 38113
rect 294811 38085 298248 38113
rect 298276 38085 298310 38113
rect 298338 38085 298372 38113
rect 298400 38085 298434 38113
rect 298462 38085 298990 38113
rect -958 38051 298990 38085
rect -958 38023 -430 38051
rect -402 38023 -368 38051
rect -340 38023 -306 38051
rect -278 38023 -244 38051
rect -216 38023 2757 38051
rect 2785 38023 2819 38051
rect 2847 38023 2881 38051
rect 2909 38023 2943 38051
rect 2971 38023 18117 38051
rect 18145 38023 18179 38051
rect 18207 38023 18241 38051
rect 18269 38023 18303 38051
rect 18331 38023 33477 38051
rect 33505 38023 33539 38051
rect 33567 38023 33601 38051
rect 33629 38023 33663 38051
rect 33691 38023 48837 38051
rect 48865 38023 48899 38051
rect 48927 38023 48961 38051
rect 48989 38023 49023 38051
rect 49051 38023 64197 38051
rect 64225 38023 64259 38051
rect 64287 38023 64321 38051
rect 64349 38023 64383 38051
rect 64411 38023 79557 38051
rect 79585 38023 79619 38051
rect 79647 38023 79681 38051
rect 79709 38023 79743 38051
rect 79771 38023 94917 38051
rect 94945 38023 94979 38051
rect 95007 38023 95041 38051
rect 95069 38023 95103 38051
rect 95131 38023 110277 38051
rect 110305 38023 110339 38051
rect 110367 38023 110401 38051
rect 110429 38023 110463 38051
rect 110491 38023 125637 38051
rect 125665 38023 125699 38051
rect 125727 38023 125761 38051
rect 125789 38023 125823 38051
rect 125851 38023 140997 38051
rect 141025 38023 141059 38051
rect 141087 38023 141121 38051
rect 141149 38023 141183 38051
rect 141211 38023 156357 38051
rect 156385 38023 156419 38051
rect 156447 38023 156481 38051
rect 156509 38023 156543 38051
rect 156571 38023 162259 38051
rect 162287 38023 162321 38051
rect 162349 38023 177619 38051
rect 177647 38023 177681 38051
rect 177709 38023 192979 38051
rect 193007 38023 193041 38051
rect 193069 38023 208339 38051
rect 208367 38023 208401 38051
rect 208429 38023 223699 38051
rect 223727 38023 223761 38051
rect 223789 38023 239059 38051
rect 239087 38023 239121 38051
rect 239149 38023 254419 38051
rect 254447 38023 254481 38051
rect 254509 38023 269779 38051
rect 269807 38023 269841 38051
rect 269869 38023 279237 38051
rect 279265 38023 279299 38051
rect 279327 38023 279361 38051
rect 279389 38023 279423 38051
rect 279451 38023 294597 38051
rect 294625 38023 294659 38051
rect 294687 38023 294721 38051
rect 294749 38023 294783 38051
rect 294811 38023 298248 38051
rect 298276 38023 298310 38051
rect 298338 38023 298372 38051
rect 298400 38023 298434 38051
rect 298462 38023 298990 38051
rect -958 37989 298990 38023
rect -958 37961 -430 37989
rect -402 37961 -368 37989
rect -340 37961 -306 37989
rect -278 37961 -244 37989
rect -216 37961 2757 37989
rect 2785 37961 2819 37989
rect 2847 37961 2881 37989
rect 2909 37961 2943 37989
rect 2971 37961 18117 37989
rect 18145 37961 18179 37989
rect 18207 37961 18241 37989
rect 18269 37961 18303 37989
rect 18331 37961 33477 37989
rect 33505 37961 33539 37989
rect 33567 37961 33601 37989
rect 33629 37961 33663 37989
rect 33691 37961 48837 37989
rect 48865 37961 48899 37989
rect 48927 37961 48961 37989
rect 48989 37961 49023 37989
rect 49051 37961 64197 37989
rect 64225 37961 64259 37989
rect 64287 37961 64321 37989
rect 64349 37961 64383 37989
rect 64411 37961 79557 37989
rect 79585 37961 79619 37989
rect 79647 37961 79681 37989
rect 79709 37961 79743 37989
rect 79771 37961 94917 37989
rect 94945 37961 94979 37989
rect 95007 37961 95041 37989
rect 95069 37961 95103 37989
rect 95131 37961 110277 37989
rect 110305 37961 110339 37989
rect 110367 37961 110401 37989
rect 110429 37961 110463 37989
rect 110491 37961 125637 37989
rect 125665 37961 125699 37989
rect 125727 37961 125761 37989
rect 125789 37961 125823 37989
rect 125851 37961 140997 37989
rect 141025 37961 141059 37989
rect 141087 37961 141121 37989
rect 141149 37961 141183 37989
rect 141211 37961 156357 37989
rect 156385 37961 156419 37989
rect 156447 37961 156481 37989
rect 156509 37961 156543 37989
rect 156571 37961 162259 37989
rect 162287 37961 162321 37989
rect 162349 37961 177619 37989
rect 177647 37961 177681 37989
rect 177709 37961 192979 37989
rect 193007 37961 193041 37989
rect 193069 37961 208339 37989
rect 208367 37961 208401 37989
rect 208429 37961 223699 37989
rect 223727 37961 223761 37989
rect 223789 37961 239059 37989
rect 239087 37961 239121 37989
rect 239149 37961 254419 37989
rect 254447 37961 254481 37989
rect 254509 37961 269779 37989
rect 269807 37961 269841 37989
rect 269869 37961 279237 37989
rect 279265 37961 279299 37989
rect 279327 37961 279361 37989
rect 279389 37961 279423 37989
rect 279451 37961 294597 37989
rect 294625 37961 294659 37989
rect 294687 37961 294721 37989
rect 294749 37961 294783 37989
rect 294811 37961 298248 37989
rect 298276 37961 298310 37989
rect 298338 37961 298372 37989
rect 298400 37961 298434 37989
rect 298462 37961 298990 37989
rect -958 37913 298990 37961
rect -958 32175 298990 32223
rect -958 32147 -910 32175
rect -882 32147 -848 32175
rect -820 32147 -786 32175
rect -758 32147 -724 32175
rect -696 32147 4617 32175
rect 4645 32147 4679 32175
rect 4707 32147 4741 32175
rect 4769 32147 4803 32175
rect 4831 32147 19977 32175
rect 20005 32147 20039 32175
rect 20067 32147 20101 32175
rect 20129 32147 20163 32175
rect 20191 32147 35337 32175
rect 35365 32147 35399 32175
rect 35427 32147 35461 32175
rect 35489 32147 35523 32175
rect 35551 32147 50697 32175
rect 50725 32147 50759 32175
rect 50787 32147 50821 32175
rect 50849 32147 50883 32175
rect 50911 32147 66057 32175
rect 66085 32147 66119 32175
rect 66147 32147 66181 32175
rect 66209 32147 66243 32175
rect 66271 32147 81417 32175
rect 81445 32147 81479 32175
rect 81507 32147 81541 32175
rect 81569 32147 81603 32175
rect 81631 32147 96777 32175
rect 96805 32147 96839 32175
rect 96867 32147 96901 32175
rect 96929 32147 96963 32175
rect 96991 32147 112137 32175
rect 112165 32147 112199 32175
rect 112227 32147 112261 32175
rect 112289 32147 112323 32175
rect 112351 32147 127497 32175
rect 127525 32147 127559 32175
rect 127587 32147 127621 32175
rect 127649 32147 127683 32175
rect 127711 32147 142857 32175
rect 142885 32147 142919 32175
rect 142947 32147 142981 32175
rect 143009 32147 143043 32175
rect 143071 32147 158217 32175
rect 158245 32147 158279 32175
rect 158307 32147 158341 32175
rect 158369 32147 158403 32175
rect 158431 32147 169939 32175
rect 169967 32147 170001 32175
rect 170029 32147 185299 32175
rect 185327 32147 185361 32175
rect 185389 32147 200659 32175
rect 200687 32147 200721 32175
rect 200749 32147 216019 32175
rect 216047 32147 216081 32175
rect 216109 32147 231379 32175
rect 231407 32147 231441 32175
rect 231469 32147 246739 32175
rect 246767 32147 246801 32175
rect 246829 32147 262099 32175
rect 262127 32147 262161 32175
rect 262189 32147 281097 32175
rect 281125 32147 281159 32175
rect 281187 32147 281221 32175
rect 281249 32147 281283 32175
rect 281311 32147 296457 32175
rect 296485 32147 296519 32175
rect 296547 32147 296581 32175
rect 296609 32147 296643 32175
rect 296671 32147 298728 32175
rect 298756 32147 298790 32175
rect 298818 32147 298852 32175
rect 298880 32147 298914 32175
rect 298942 32147 298990 32175
rect -958 32113 298990 32147
rect -958 32085 -910 32113
rect -882 32085 -848 32113
rect -820 32085 -786 32113
rect -758 32085 -724 32113
rect -696 32085 4617 32113
rect 4645 32085 4679 32113
rect 4707 32085 4741 32113
rect 4769 32085 4803 32113
rect 4831 32085 19977 32113
rect 20005 32085 20039 32113
rect 20067 32085 20101 32113
rect 20129 32085 20163 32113
rect 20191 32085 35337 32113
rect 35365 32085 35399 32113
rect 35427 32085 35461 32113
rect 35489 32085 35523 32113
rect 35551 32085 50697 32113
rect 50725 32085 50759 32113
rect 50787 32085 50821 32113
rect 50849 32085 50883 32113
rect 50911 32085 66057 32113
rect 66085 32085 66119 32113
rect 66147 32085 66181 32113
rect 66209 32085 66243 32113
rect 66271 32085 81417 32113
rect 81445 32085 81479 32113
rect 81507 32085 81541 32113
rect 81569 32085 81603 32113
rect 81631 32085 96777 32113
rect 96805 32085 96839 32113
rect 96867 32085 96901 32113
rect 96929 32085 96963 32113
rect 96991 32085 112137 32113
rect 112165 32085 112199 32113
rect 112227 32085 112261 32113
rect 112289 32085 112323 32113
rect 112351 32085 127497 32113
rect 127525 32085 127559 32113
rect 127587 32085 127621 32113
rect 127649 32085 127683 32113
rect 127711 32085 142857 32113
rect 142885 32085 142919 32113
rect 142947 32085 142981 32113
rect 143009 32085 143043 32113
rect 143071 32085 158217 32113
rect 158245 32085 158279 32113
rect 158307 32085 158341 32113
rect 158369 32085 158403 32113
rect 158431 32085 169939 32113
rect 169967 32085 170001 32113
rect 170029 32085 185299 32113
rect 185327 32085 185361 32113
rect 185389 32085 200659 32113
rect 200687 32085 200721 32113
rect 200749 32085 216019 32113
rect 216047 32085 216081 32113
rect 216109 32085 231379 32113
rect 231407 32085 231441 32113
rect 231469 32085 246739 32113
rect 246767 32085 246801 32113
rect 246829 32085 262099 32113
rect 262127 32085 262161 32113
rect 262189 32085 281097 32113
rect 281125 32085 281159 32113
rect 281187 32085 281221 32113
rect 281249 32085 281283 32113
rect 281311 32085 296457 32113
rect 296485 32085 296519 32113
rect 296547 32085 296581 32113
rect 296609 32085 296643 32113
rect 296671 32085 298728 32113
rect 298756 32085 298790 32113
rect 298818 32085 298852 32113
rect 298880 32085 298914 32113
rect 298942 32085 298990 32113
rect -958 32051 298990 32085
rect -958 32023 -910 32051
rect -882 32023 -848 32051
rect -820 32023 -786 32051
rect -758 32023 -724 32051
rect -696 32023 4617 32051
rect 4645 32023 4679 32051
rect 4707 32023 4741 32051
rect 4769 32023 4803 32051
rect 4831 32023 19977 32051
rect 20005 32023 20039 32051
rect 20067 32023 20101 32051
rect 20129 32023 20163 32051
rect 20191 32023 35337 32051
rect 35365 32023 35399 32051
rect 35427 32023 35461 32051
rect 35489 32023 35523 32051
rect 35551 32023 50697 32051
rect 50725 32023 50759 32051
rect 50787 32023 50821 32051
rect 50849 32023 50883 32051
rect 50911 32023 66057 32051
rect 66085 32023 66119 32051
rect 66147 32023 66181 32051
rect 66209 32023 66243 32051
rect 66271 32023 81417 32051
rect 81445 32023 81479 32051
rect 81507 32023 81541 32051
rect 81569 32023 81603 32051
rect 81631 32023 96777 32051
rect 96805 32023 96839 32051
rect 96867 32023 96901 32051
rect 96929 32023 96963 32051
rect 96991 32023 112137 32051
rect 112165 32023 112199 32051
rect 112227 32023 112261 32051
rect 112289 32023 112323 32051
rect 112351 32023 127497 32051
rect 127525 32023 127559 32051
rect 127587 32023 127621 32051
rect 127649 32023 127683 32051
rect 127711 32023 142857 32051
rect 142885 32023 142919 32051
rect 142947 32023 142981 32051
rect 143009 32023 143043 32051
rect 143071 32023 158217 32051
rect 158245 32023 158279 32051
rect 158307 32023 158341 32051
rect 158369 32023 158403 32051
rect 158431 32023 169939 32051
rect 169967 32023 170001 32051
rect 170029 32023 185299 32051
rect 185327 32023 185361 32051
rect 185389 32023 200659 32051
rect 200687 32023 200721 32051
rect 200749 32023 216019 32051
rect 216047 32023 216081 32051
rect 216109 32023 231379 32051
rect 231407 32023 231441 32051
rect 231469 32023 246739 32051
rect 246767 32023 246801 32051
rect 246829 32023 262099 32051
rect 262127 32023 262161 32051
rect 262189 32023 281097 32051
rect 281125 32023 281159 32051
rect 281187 32023 281221 32051
rect 281249 32023 281283 32051
rect 281311 32023 296457 32051
rect 296485 32023 296519 32051
rect 296547 32023 296581 32051
rect 296609 32023 296643 32051
rect 296671 32023 298728 32051
rect 298756 32023 298790 32051
rect 298818 32023 298852 32051
rect 298880 32023 298914 32051
rect 298942 32023 298990 32051
rect -958 31989 298990 32023
rect -958 31961 -910 31989
rect -882 31961 -848 31989
rect -820 31961 -786 31989
rect -758 31961 -724 31989
rect -696 31961 4617 31989
rect 4645 31961 4679 31989
rect 4707 31961 4741 31989
rect 4769 31961 4803 31989
rect 4831 31961 19977 31989
rect 20005 31961 20039 31989
rect 20067 31961 20101 31989
rect 20129 31961 20163 31989
rect 20191 31961 35337 31989
rect 35365 31961 35399 31989
rect 35427 31961 35461 31989
rect 35489 31961 35523 31989
rect 35551 31961 50697 31989
rect 50725 31961 50759 31989
rect 50787 31961 50821 31989
rect 50849 31961 50883 31989
rect 50911 31961 66057 31989
rect 66085 31961 66119 31989
rect 66147 31961 66181 31989
rect 66209 31961 66243 31989
rect 66271 31961 81417 31989
rect 81445 31961 81479 31989
rect 81507 31961 81541 31989
rect 81569 31961 81603 31989
rect 81631 31961 96777 31989
rect 96805 31961 96839 31989
rect 96867 31961 96901 31989
rect 96929 31961 96963 31989
rect 96991 31961 112137 31989
rect 112165 31961 112199 31989
rect 112227 31961 112261 31989
rect 112289 31961 112323 31989
rect 112351 31961 127497 31989
rect 127525 31961 127559 31989
rect 127587 31961 127621 31989
rect 127649 31961 127683 31989
rect 127711 31961 142857 31989
rect 142885 31961 142919 31989
rect 142947 31961 142981 31989
rect 143009 31961 143043 31989
rect 143071 31961 158217 31989
rect 158245 31961 158279 31989
rect 158307 31961 158341 31989
rect 158369 31961 158403 31989
rect 158431 31961 169939 31989
rect 169967 31961 170001 31989
rect 170029 31961 185299 31989
rect 185327 31961 185361 31989
rect 185389 31961 200659 31989
rect 200687 31961 200721 31989
rect 200749 31961 216019 31989
rect 216047 31961 216081 31989
rect 216109 31961 231379 31989
rect 231407 31961 231441 31989
rect 231469 31961 246739 31989
rect 246767 31961 246801 31989
rect 246829 31961 262099 31989
rect 262127 31961 262161 31989
rect 262189 31961 281097 31989
rect 281125 31961 281159 31989
rect 281187 31961 281221 31989
rect 281249 31961 281283 31989
rect 281311 31961 296457 31989
rect 296485 31961 296519 31989
rect 296547 31961 296581 31989
rect 296609 31961 296643 31989
rect 296671 31961 298728 31989
rect 298756 31961 298790 31989
rect 298818 31961 298852 31989
rect 298880 31961 298914 31989
rect 298942 31961 298990 31989
rect -958 31913 298990 31961
rect -958 29175 298990 29223
rect -958 29147 -430 29175
rect -402 29147 -368 29175
rect -340 29147 -306 29175
rect -278 29147 -244 29175
rect -216 29147 2757 29175
rect 2785 29147 2819 29175
rect 2847 29147 2881 29175
rect 2909 29147 2943 29175
rect 2971 29147 18117 29175
rect 18145 29147 18179 29175
rect 18207 29147 18241 29175
rect 18269 29147 18303 29175
rect 18331 29147 33477 29175
rect 33505 29147 33539 29175
rect 33567 29147 33601 29175
rect 33629 29147 33663 29175
rect 33691 29147 48837 29175
rect 48865 29147 48899 29175
rect 48927 29147 48961 29175
rect 48989 29147 49023 29175
rect 49051 29147 64197 29175
rect 64225 29147 64259 29175
rect 64287 29147 64321 29175
rect 64349 29147 64383 29175
rect 64411 29147 79557 29175
rect 79585 29147 79619 29175
rect 79647 29147 79681 29175
rect 79709 29147 79743 29175
rect 79771 29147 94917 29175
rect 94945 29147 94979 29175
rect 95007 29147 95041 29175
rect 95069 29147 95103 29175
rect 95131 29147 110277 29175
rect 110305 29147 110339 29175
rect 110367 29147 110401 29175
rect 110429 29147 110463 29175
rect 110491 29147 125637 29175
rect 125665 29147 125699 29175
rect 125727 29147 125761 29175
rect 125789 29147 125823 29175
rect 125851 29147 140997 29175
rect 141025 29147 141059 29175
rect 141087 29147 141121 29175
rect 141149 29147 141183 29175
rect 141211 29147 156357 29175
rect 156385 29147 156419 29175
rect 156447 29147 156481 29175
rect 156509 29147 156543 29175
rect 156571 29147 162259 29175
rect 162287 29147 162321 29175
rect 162349 29147 177619 29175
rect 177647 29147 177681 29175
rect 177709 29147 192979 29175
rect 193007 29147 193041 29175
rect 193069 29147 208339 29175
rect 208367 29147 208401 29175
rect 208429 29147 223699 29175
rect 223727 29147 223761 29175
rect 223789 29147 239059 29175
rect 239087 29147 239121 29175
rect 239149 29147 254419 29175
rect 254447 29147 254481 29175
rect 254509 29147 269779 29175
rect 269807 29147 269841 29175
rect 269869 29147 279237 29175
rect 279265 29147 279299 29175
rect 279327 29147 279361 29175
rect 279389 29147 279423 29175
rect 279451 29147 294597 29175
rect 294625 29147 294659 29175
rect 294687 29147 294721 29175
rect 294749 29147 294783 29175
rect 294811 29147 298248 29175
rect 298276 29147 298310 29175
rect 298338 29147 298372 29175
rect 298400 29147 298434 29175
rect 298462 29147 298990 29175
rect -958 29113 298990 29147
rect -958 29085 -430 29113
rect -402 29085 -368 29113
rect -340 29085 -306 29113
rect -278 29085 -244 29113
rect -216 29085 2757 29113
rect 2785 29085 2819 29113
rect 2847 29085 2881 29113
rect 2909 29085 2943 29113
rect 2971 29085 18117 29113
rect 18145 29085 18179 29113
rect 18207 29085 18241 29113
rect 18269 29085 18303 29113
rect 18331 29085 33477 29113
rect 33505 29085 33539 29113
rect 33567 29085 33601 29113
rect 33629 29085 33663 29113
rect 33691 29085 48837 29113
rect 48865 29085 48899 29113
rect 48927 29085 48961 29113
rect 48989 29085 49023 29113
rect 49051 29085 64197 29113
rect 64225 29085 64259 29113
rect 64287 29085 64321 29113
rect 64349 29085 64383 29113
rect 64411 29085 79557 29113
rect 79585 29085 79619 29113
rect 79647 29085 79681 29113
rect 79709 29085 79743 29113
rect 79771 29085 94917 29113
rect 94945 29085 94979 29113
rect 95007 29085 95041 29113
rect 95069 29085 95103 29113
rect 95131 29085 110277 29113
rect 110305 29085 110339 29113
rect 110367 29085 110401 29113
rect 110429 29085 110463 29113
rect 110491 29085 125637 29113
rect 125665 29085 125699 29113
rect 125727 29085 125761 29113
rect 125789 29085 125823 29113
rect 125851 29085 140997 29113
rect 141025 29085 141059 29113
rect 141087 29085 141121 29113
rect 141149 29085 141183 29113
rect 141211 29085 156357 29113
rect 156385 29085 156419 29113
rect 156447 29085 156481 29113
rect 156509 29085 156543 29113
rect 156571 29085 162259 29113
rect 162287 29085 162321 29113
rect 162349 29085 177619 29113
rect 177647 29085 177681 29113
rect 177709 29085 192979 29113
rect 193007 29085 193041 29113
rect 193069 29085 208339 29113
rect 208367 29085 208401 29113
rect 208429 29085 223699 29113
rect 223727 29085 223761 29113
rect 223789 29085 239059 29113
rect 239087 29085 239121 29113
rect 239149 29085 254419 29113
rect 254447 29085 254481 29113
rect 254509 29085 269779 29113
rect 269807 29085 269841 29113
rect 269869 29085 279237 29113
rect 279265 29085 279299 29113
rect 279327 29085 279361 29113
rect 279389 29085 279423 29113
rect 279451 29085 294597 29113
rect 294625 29085 294659 29113
rect 294687 29085 294721 29113
rect 294749 29085 294783 29113
rect 294811 29085 298248 29113
rect 298276 29085 298310 29113
rect 298338 29085 298372 29113
rect 298400 29085 298434 29113
rect 298462 29085 298990 29113
rect -958 29051 298990 29085
rect -958 29023 -430 29051
rect -402 29023 -368 29051
rect -340 29023 -306 29051
rect -278 29023 -244 29051
rect -216 29023 2757 29051
rect 2785 29023 2819 29051
rect 2847 29023 2881 29051
rect 2909 29023 2943 29051
rect 2971 29023 18117 29051
rect 18145 29023 18179 29051
rect 18207 29023 18241 29051
rect 18269 29023 18303 29051
rect 18331 29023 33477 29051
rect 33505 29023 33539 29051
rect 33567 29023 33601 29051
rect 33629 29023 33663 29051
rect 33691 29023 48837 29051
rect 48865 29023 48899 29051
rect 48927 29023 48961 29051
rect 48989 29023 49023 29051
rect 49051 29023 64197 29051
rect 64225 29023 64259 29051
rect 64287 29023 64321 29051
rect 64349 29023 64383 29051
rect 64411 29023 79557 29051
rect 79585 29023 79619 29051
rect 79647 29023 79681 29051
rect 79709 29023 79743 29051
rect 79771 29023 94917 29051
rect 94945 29023 94979 29051
rect 95007 29023 95041 29051
rect 95069 29023 95103 29051
rect 95131 29023 110277 29051
rect 110305 29023 110339 29051
rect 110367 29023 110401 29051
rect 110429 29023 110463 29051
rect 110491 29023 125637 29051
rect 125665 29023 125699 29051
rect 125727 29023 125761 29051
rect 125789 29023 125823 29051
rect 125851 29023 140997 29051
rect 141025 29023 141059 29051
rect 141087 29023 141121 29051
rect 141149 29023 141183 29051
rect 141211 29023 156357 29051
rect 156385 29023 156419 29051
rect 156447 29023 156481 29051
rect 156509 29023 156543 29051
rect 156571 29023 162259 29051
rect 162287 29023 162321 29051
rect 162349 29023 177619 29051
rect 177647 29023 177681 29051
rect 177709 29023 192979 29051
rect 193007 29023 193041 29051
rect 193069 29023 208339 29051
rect 208367 29023 208401 29051
rect 208429 29023 223699 29051
rect 223727 29023 223761 29051
rect 223789 29023 239059 29051
rect 239087 29023 239121 29051
rect 239149 29023 254419 29051
rect 254447 29023 254481 29051
rect 254509 29023 269779 29051
rect 269807 29023 269841 29051
rect 269869 29023 279237 29051
rect 279265 29023 279299 29051
rect 279327 29023 279361 29051
rect 279389 29023 279423 29051
rect 279451 29023 294597 29051
rect 294625 29023 294659 29051
rect 294687 29023 294721 29051
rect 294749 29023 294783 29051
rect 294811 29023 298248 29051
rect 298276 29023 298310 29051
rect 298338 29023 298372 29051
rect 298400 29023 298434 29051
rect 298462 29023 298990 29051
rect -958 28989 298990 29023
rect -958 28961 -430 28989
rect -402 28961 -368 28989
rect -340 28961 -306 28989
rect -278 28961 -244 28989
rect -216 28961 2757 28989
rect 2785 28961 2819 28989
rect 2847 28961 2881 28989
rect 2909 28961 2943 28989
rect 2971 28961 18117 28989
rect 18145 28961 18179 28989
rect 18207 28961 18241 28989
rect 18269 28961 18303 28989
rect 18331 28961 33477 28989
rect 33505 28961 33539 28989
rect 33567 28961 33601 28989
rect 33629 28961 33663 28989
rect 33691 28961 48837 28989
rect 48865 28961 48899 28989
rect 48927 28961 48961 28989
rect 48989 28961 49023 28989
rect 49051 28961 64197 28989
rect 64225 28961 64259 28989
rect 64287 28961 64321 28989
rect 64349 28961 64383 28989
rect 64411 28961 79557 28989
rect 79585 28961 79619 28989
rect 79647 28961 79681 28989
rect 79709 28961 79743 28989
rect 79771 28961 94917 28989
rect 94945 28961 94979 28989
rect 95007 28961 95041 28989
rect 95069 28961 95103 28989
rect 95131 28961 110277 28989
rect 110305 28961 110339 28989
rect 110367 28961 110401 28989
rect 110429 28961 110463 28989
rect 110491 28961 125637 28989
rect 125665 28961 125699 28989
rect 125727 28961 125761 28989
rect 125789 28961 125823 28989
rect 125851 28961 140997 28989
rect 141025 28961 141059 28989
rect 141087 28961 141121 28989
rect 141149 28961 141183 28989
rect 141211 28961 156357 28989
rect 156385 28961 156419 28989
rect 156447 28961 156481 28989
rect 156509 28961 156543 28989
rect 156571 28961 162259 28989
rect 162287 28961 162321 28989
rect 162349 28961 177619 28989
rect 177647 28961 177681 28989
rect 177709 28961 192979 28989
rect 193007 28961 193041 28989
rect 193069 28961 208339 28989
rect 208367 28961 208401 28989
rect 208429 28961 223699 28989
rect 223727 28961 223761 28989
rect 223789 28961 239059 28989
rect 239087 28961 239121 28989
rect 239149 28961 254419 28989
rect 254447 28961 254481 28989
rect 254509 28961 269779 28989
rect 269807 28961 269841 28989
rect 269869 28961 279237 28989
rect 279265 28961 279299 28989
rect 279327 28961 279361 28989
rect 279389 28961 279423 28989
rect 279451 28961 294597 28989
rect 294625 28961 294659 28989
rect 294687 28961 294721 28989
rect 294749 28961 294783 28989
rect 294811 28961 298248 28989
rect 298276 28961 298310 28989
rect 298338 28961 298372 28989
rect 298400 28961 298434 28989
rect 298462 28961 298990 28989
rect -958 28913 298990 28961
rect -958 23175 298990 23223
rect -958 23147 -910 23175
rect -882 23147 -848 23175
rect -820 23147 -786 23175
rect -758 23147 -724 23175
rect -696 23147 4617 23175
rect 4645 23147 4679 23175
rect 4707 23147 4741 23175
rect 4769 23147 4803 23175
rect 4831 23147 19977 23175
rect 20005 23147 20039 23175
rect 20067 23147 20101 23175
rect 20129 23147 20163 23175
rect 20191 23147 35337 23175
rect 35365 23147 35399 23175
rect 35427 23147 35461 23175
rect 35489 23147 35523 23175
rect 35551 23147 50697 23175
rect 50725 23147 50759 23175
rect 50787 23147 50821 23175
rect 50849 23147 50883 23175
rect 50911 23147 66057 23175
rect 66085 23147 66119 23175
rect 66147 23147 66181 23175
rect 66209 23147 66243 23175
rect 66271 23147 81417 23175
rect 81445 23147 81479 23175
rect 81507 23147 81541 23175
rect 81569 23147 81603 23175
rect 81631 23147 96777 23175
rect 96805 23147 96839 23175
rect 96867 23147 96901 23175
rect 96929 23147 96963 23175
rect 96991 23147 112137 23175
rect 112165 23147 112199 23175
rect 112227 23147 112261 23175
rect 112289 23147 112323 23175
rect 112351 23147 127497 23175
rect 127525 23147 127559 23175
rect 127587 23147 127621 23175
rect 127649 23147 127683 23175
rect 127711 23147 142857 23175
rect 142885 23147 142919 23175
rect 142947 23147 142981 23175
rect 143009 23147 143043 23175
rect 143071 23147 158217 23175
rect 158245 23147 158279 23175
rect 158307 23147 158341 23175
rect 158369 23147 158403 23175
rect 158431 23147 169939 23175
rect 169967 23147 170001 23175
rect 170029 23147 185299 23175
rect 185327 23147 185361 23175
rect 185389 23147 200659 23175
rect 200687 23147 200721 23175
rect 200749 23147 216019 23175
rect 216047 23147 216081 23175
rect 216109 23147 231379 23175
rect 231407 23147 231441 23175
rect 231469 23147 246739 23175
rect 246767 23147 246801 23175
rect 246829 23147 262099 23175
rect 262127 23147 262161 23175
rect 262189 23147 281097 23175
rect 281125 23147 281159 23175
rect 281187 23147 281221 23175
rect 281249 23147 281283 23175
rect 281311 23147 296457 23175
rect 296485 23147 296519 23175
rect 296547 23147 296581 23175
rect 296609 23147 296643 23175
rect 296671 23147 298728 23175
rect 298756 23147 298790 23175
rect 298818 23147 298852 23175
rect 298880 23147 298914 23175
rect 298942 23147 298990 23175
rect -958 23113 298990 23147
rect -958 23085 -910 23113
rect -882 23085 -848 23113
rect -820 23085 -786 23113
rect -758 23085 -724 23113
rect -696 23085 4617 23113
rect 4645 23085 4679 23113
rect 4707 23085 4741 23113
rect 4769 23085 4803 23113
rect 4831 23085 19977 23113
rect 20005 23085 20039 23113
rect 20067 23085 20101 23113
rect 20129 23085 20163 23113
rect 20191 23085 35337 23113
rect 35365 23085 35399 23113
rect 35427 23085 35461 23113
rect 35489 23085 35523 23113
rect 35551 23085 50697 23113
rect 50725 23085 50759 23113
rect 50787 23085 50821 23113
rect 50849 23085 50883 23113
rect 50911 23085 66057 23113
rect 66085 23085 66119 23113
rect 66147 23085 66181 23113
rect 66209 23085 66243 23113
rect 66271 23085 81417 23113
rect 81445 23085 81479 23113
rect 81507 23085 81541 23113
rect 81569 23085 81603 23113
rect 81631 23085 96777 23113
rect 96805 23085 96839 23113
rect 96867 23085 96901 23113
rect 96929 23085 96963 23113
rect 96991 23085 112137 23113
rect 112165 23085 112199 23113
rect 112227 23085 112261 23113
rect 112289 23085 112323 23113
rect 112351 23085 127497 23113
rect 127525 23085 127559 23113
rect 127587 23085 127621 23113
rect 127649 23085 127683 23113
rect 127711 23085 142857 23113
rect 142885 23085 142919 23113
rect 142947 23085 142981 23113
rect 143009 23085 143043 23113
rect 143071 23085 158217 23113
rect 158245 23085 158279 23113
rect 158307 23085 158341 23113
rect 158369 23085 158403 23113
rect 158431 23085 169939 23113
rect 169967 23085 170001 23113
rect 170029 23085 185299 23113
rect 185327 23085 185361 23113
rect 185389 23085 200659 23113
rect 200687 23085 200721 23113
rect 200749 23085 216019 23113
rect 216047 23085 216081 23113
rect 216109 23085 231379 23113
rect 231407 23085 231441 23113
rect 231469 23085 246739 23113
rect 246767 23085 246801 23113
rect 246829 23085 262099 23113
rect 262127 23085 262161 23113
rect 262189 23085 281097 23113
rect 281125 23085 281159 23113
rect 281187 23085 281221 23113
rect 281249 23085 281283 23113
rect 281311 23085 296457 23113
rect 296485 23085 296519 23113
rect 296547 23085 296581 23113
rect 296609 23085 296643 23113
rect 296671 23085 298728 23113
rect 298756 23085 298790 23113
rect 298818 23085 298852 23113
rect 298880 23085 298914 23113
rect 298942 23085 298990 23113
rect -958 23051 298990 23085
rect -958 23023 -910 23051
rect -882 23023 -848 23051
rect -820 23023 -786 23051
rect -758 23023 -724 23051
rect -696 23023 4617 23051
rect 4645 23023 4679 23051
rect 4707 23023 4741 23051
rect 4769 23023 4803 23051
rect 4831 23023 19977 23051
rect 20005 23023 20039 23051
rect 20067 23023 20101 23051
rect 20129 23023 20163 23051
rect 20191 23023 35337 23051
rect 35365 23023 35399 23051
rect 35427 23023 35461 23051
rect 35489 23023 35523 23051
rect 35551 23023 50697 23051
rect 50725 23023 50759 23051
rect 50787 23023 50821 23051
rect 50849 23023 50883 23051
rect 50911 23023 66057 23051
rect 66085 23023 66119 23051
rect 66147 23023 66181 23051
rect 66209 23023 66243 23051
rect 66271 23023 81417 23051
rect 81445 23023 81479 23051
rect 81507 23023 81541 23051
rect 81569 23023 81603 23051
rect 81631 23023 96777 23051
rect 96805 23023 96839 23051
rect 96867 23023 96901 23051
rect 96929 23023 96963 23051
rect 96991 23023 112137 23051
rect 112165 23023 112199 23051
rect 112227 23023 112261 23051
rect 112289 23023 112323 23051
rect 112351 23023 127497 23051
rect 127525 23023 127559 23051
rect 127587 23023 127621 23051
rect 127649 23023 127683 23051
rect 127711 23023 142857 23051
rect 142885 23023 142919 23051
rect 142947 23023 142981 23051
rect 143009 23023 143043 23051
rect 143071 23023 158217 23051
rect 158245 23023 158279 23051
rect 158307 23023 158341 23051
rect 158369 23023 158403 23051
rect 158431 23023 169939 23051
rect 169967 23023 170001 23051
rect 170029 23023 185299 23051
rect 185327 23023 185361 23051
rect 185389 23023 200659 23051
rect 200687 23023 200721 23051
rect 200749 23023 216019 23051
rect 216047 23023 216081 23051
rect 216109 23023 231379 23051
rect 231407 23023 231441 23051
rect 231469 23023 246739 23051
rect 246767 23023 246801 23051
rect 246829 23023 262099 23051
rect 262127 23023 262161 23051
rect 262189 23023 281097 23051
rect 281125 23023 281159 23051
rect 281187 23023 281221 23051
rect 281249 23023 281283 23051
rect 281311 23023 296457 23051
rect 296485 23023 296519 23051
rect 296547 23023 296581 23051
rect 296609 23023 296643 23051
rect 296671 23023 298728 23051
rect 298756 23023 298790 23051
rect 298818 23023 298852 23051
rect 298880 23023 298914 23051
rect 298942 23023 298990 23051
rect -958 22989 298990 23023
rect -958 22961 -910 22989
rect -882 22961 -848 22989
rect -820 22961 -786 22989
rect -758 22961 -724 22989
rect -696 22961 4617 22989
rect 4645 22961 4679 22989
rect 4707 22961 4741 22989
rect 4769 22961 4803 22989
rect 4831 22961 19977 22989
rect 20005 22961 20039 22989
rect 20067 22961 20101 22989
rect 20129 22961 20163 22989
rect 20191 22961 35337 22989
rect 35365 22961 35399 22989
rect 35427 22961 35461 22989
rect 35489 22961 35523 22989
rect 35551 22961 50697 22989
rect 50725 22961 50759 22989
rect 50787 22961 50821 22989
rect 50849 22961 50883 22989
rect 50911 22961 66057 22989
rect 66085 22961 66119 22989
rect 66147 22961 66181 22989
rect 66209 22961 66243 22989
rect 66271 22961 81417 22989
rect 81445 22961 81479 22989
rect 81507 22961 81541 22989
rect 81569 22961 81603 22989
rect 81631 22961 96777 22989
rect 96805 22961 96839 22989
rect 96867 22961 96901 22989
rect 96929 22961 96963 22989
rect 96991 22961 112137 22989
rect 112165 22961 112199 22989
rect 112227 22961 112261 22989
rect 112289 22961 112323 22989
rect 112351 22961 127497 22989
rect 127525 22961 127559 22989
rect 127587 22961 127621 22989
rect 127649 22961 127683 22989
rect 127711 22961 142857 22989
rect 142885 22961 142919 22989
rect 142947 22961 142981 22989
rect 143009 22961 143043 22989
rect 143071 22961 158217 22989
rect 158245 22961 158279 22989
rect 158307 22961 158341 22989
rect 158369 22961 158403 22989
rect 158431 22961 169939 22989
rect 169967 22961 170001 22989
rect 170029 22961 185299 22989
rect 185327 22961 185361 22989
rect 185389 22961 200659 22989
rect 200687 22961 200721 22989
rect 200749 22961 216019 22989
rect 216047 22961 216081 22989
rect 216109 22961 231379 22989
rect 231407 22961 231441 22989
rect 231469 22961 246739 22989
rect 246767 22961 246801 22989
rect 246829 22961 262099 22989
rect 262127 22961 262161 22989
rect 262189 22961 281097 22989
rect 281125 22961 281159 22989
rect 281187 22961 281221 22989
rect 281249 22961 281283 22989
rect 281311 22961 296457 22989
rect 296485 22961 296519 22989
rect 296547 22961 296581 22989
rect 296609 22961 296643 22989
rect 296671 22961 298728 22989
rect 298756 22961 298790 22989
rect 298818 22961 298852 22989
rect 298880 22961 298914 22989
rect 298942 22961 298990 22989
rect -958 22913 298990 22961
rect -958 20175 298990 20223
rect -958 20147 -430 20175
rect -402 20147 -368 20175
rect -340 20147 -306 20175
rect -278 20147 -244 20175
rect -216 20147 2757 20175
rect 2785 20147 2819 20175
rect 2847 20147 2881 20175
rect 2909 20147 2943 20175
rect 2971 20147 18117 20175
rect 18145 20147 18179 20175
rect 18207 20147 18241 20175
rect 18269 20147 18303 20175
rect 18331 20147 33477 20175
rect 33505 20147 33539 20175
rect 33567 20147 33601 20175
rect 33629 20147 33663 20175
rect 33691 20147 48837 20175
rect 48865 20147 48899 20175
rect 48927 20147 48961 20175
rect 48989 20147 49023 20175
rect 49051 20147 64197 20175
rect 64225 20147 64259 20175
rect 64287 20147 64321 20175
rect 64349 20147 64383 20175
rect 64411 20147 79557 20175
rect 79585 20147 79619 20175
rect 79647 20147 79681 20175
rect 79709 20147 79743 20175
rect 79771 20147 94917 20175
rect 94945 20147 94979 20175
rect 95007 20147 95041 20175
rect 95069 20147 95103 20175
rect 95131 20147 110277 20175
rect 110305 20147 110339 20175
rect 110367 20147 110401 20175
rect 110429 20147 110463 20175
rect 110491 20147 125637 20175
rect 125665 20147 125699 20175
rect 125727 20147 125761 20175
rect 125789 20147 125823 20175
rect 125851 20147 140997 20175
rect 141025 20147 141059 20175
rect 141087 20147 141121 20175
rect 141149 20147 141183 20175
rect 141211 20147 156357 20175
rect 156385 20147 156419 20175
rect 156447 20147 156481 20175
rect 156509 20147 156543 20175
rect 156571 20147 162259 20175
rect 162287 20147 162321 20175
rect 162349 20147 177619 20175
rect 177647 20147 177681 20175
rect 177709 20147 192979 20175
rect 193007 20147 193041 20175
rect 193069 20147 208339 20175
rect 208367 20147 208401 20175
rect 208429 20147 223699 20175
rect 223727 20147 223761 20175
rect 223789 20147 239059 20175
rect 239087 20147 239121 20175
rect 239149 20147 254419 20175
rect 254447 20147 254481 20175
rect 254509 20147 269779 20175
rect 269807 20147 269841 20175
rect 269869 20147 279237 20175
rect 279265 20147 279299 20175
rect 279327 20147 279361 20175
rect 279389 20147 279423 20175
rect 279451 20147 294597 20175
rect 294625 20147 294659 20175
rect 294687 20147 294721 20175
rect 294749 20147 294783 20175
rect 294811 20147 298248 20175
rect 298276 20147 298310 20175
rect 298338 20147 298372 20175
rect 298400 20147 298434 20175
rect 298462 20147 298990 20175
rect -958 20113 298990 20147
rect -958 20085 -430 20113
rect -402 20085 -368 20113
rect -340 20085 -306 20113
rect -278 20085 -244 20113
rect -216 20085 2757 20113
rect 2785 20085 2819 20113
rect 2847 20085 2881 20113
rect 2909 20085 2943 20113
rect 2971 20085 18117 20113
rect 18145 20085 18179 20113
rect 18207 20085 18241 20113
rect 18269 20085 18303 20113
rect 18331 20085 33477 20113
rect 33505 20085 33539 20113
rect 33567 20085 33601 20113
rect 33629 20085 33663 20113
rect 33691 20085 48837 20113
rect 48865 20085 48899 20113
rect 48927 20085 48961 20113
rect 48989 20085 49023 20113
rect 49051 20085 64197 20113
rect 64225 20085 64259 20113
rect 64287 20085 64321 20113
rect 64349 20085 64383 20113
rect 64411 20085 79557 20113
rect 79585 20085 79619 20113
rect 79647 20085 79681 20113
rect 79709 20085 79743 20113
rect 79771 20085 94917 20113
rect 94945 20085 94979 20113
rect 95007 20085 95041 20113
rect 95069 20085 95103 20113
rect 95131 20085 110277 20113
rect 110305 20085 110339 20113
rect 110367 20085 110401 20113
rect 110429 20085 110463 20113
rect 110491 20085 125637 20113
rect 125665 20085 125699 20113
rect 125727 20085 125761 20113
rect 125789 20085 125823 20113
rect 125851 20085 140997 20113
rect 141025 20085 141059 20113
rect 141087 20085 141121 20113
rect 141149 20085 141183 20113
rect 141211 20085 156357 20113
rect 156385 20085 156419 20113
rect 156447 20085 156481 20113
rect 156509 20085 156543 20113
rect 156571 20085 162259 20113
rect 162287 20085 162321 20113
rect 162349 20085 177619 20113
rect 177647 20085 177681 20113
rect 177709 20085 192979 20113
rect 193007 20085 193041 20113
rect 193069 20085 208339 20113
rect 208367 20085 208401 20113
rect 208429 20085 223699 20113
rect 223727 20085 223761 20113
rect 223789 20085 239059 20113
rect 239087 20085 239121 20113
rect 239149 20085 254419 20113
rect 254447 20085 254481 20113
rect 254509 20085 269779 20113
rect 269807 20085 269841 20113
rect 269869 20085 279237 20113
rect 279265 20085 279299 20113
rect 279327 20085 279361 20113
rect 279389 20085 279423 20113
rect 279451 20085 294597 20113
rect 294625 20085 294659 20113
rect 294687 20085 294721 20113
rect 294749 20085 294783 20113
rect 294811 20085 298248 20113
rect 298276 20085 298310 20113
rect 298338 20085 298372 20113
rect 298400 20085 298434 20113
rect 298462 20085 298990 20113
rect -958 20051 298990 20085
rect -958 20023 -430 20051
rect -402 20023 -368 20051
rect -340 20023 -306 20051
rect -278 20023 -244 20051
rect -216 20023 2757 20051
rect 2785 20023 2819 20051
rect 2847 20023 2881 20051
rect 2909 20023 2943 20051
rect 2971 20023 18117 20051
rect 18145 20023 18179 20051
rect 18207 20023 18241 20051
rect 18269 20023 18303 20051
rect 18331 20023 33477 20051
rect 33505 20023 33539 20051
rect 33567 20023 33601 20051
rect 33629 20023 33663 20051
rect 33691 20023 48837 20051
rect 48865 20023 48899 20051
rect 48927 20023 48961 20051
rect 48989 20023 49023 20051
rect 49051 20023 64197 20051
rect 64225 20023 64259 20051
rect 64287 20023 64321 20051
rect 64349 20023 64383 20051
rect 64411 20023 79557 20051
rect 79585 20023 79619 20051
rect 79647 20023 79681 20051
rect 79709 20023 79743 20051
rect 79771 20023 94917 20051
rect 94945 20023 94979 20051
rect 95007 20023 95041 20051
rect 95069 20023 95103 20051
rect 95131 20023 110277 20051
rect 110305 20023 110339 20051
rect 110367 20023 110401 20051
rect 110429 20023 110463 20051
rect 110491 20023 125637 20051
rect 125665 20023 125699 20051
rect 125727 20023 125761 20051
rect 125789 20023 125823 20051
rect 125851 20023 140997 20051
rect 141025 20023 141059 20051
rect 141087 20023 141121 20051
rect 141149 20023 141183 20051
rect 141211 20023 156357 20051
rect 156385 20023 156419 20051
rect 156447 20023 156481 20051
rect 156509 20023 156543 20051
rect 156571 20023 162259 20051
rect 162287 20023 162321 20051
rect 162349 20023 177619 20051
rect 177647 20023 177681 20051
rect 177709 20023 192979 20051
rect 193007 20023 193041 20051
rect 193069 20023 208339 20051
rect 208367 20023 208401 20051
rect 208429 20023 223699 20051
rect 223727 20023 223761 20051
rect 223789 20023 239059 20051
rect 239087 20023 239121 20051
rect 239149 20023 254419 20051
rect 254447 20023 254481 20051
rect 254509 20023 269779 20051
rect 269807 20023 269841 20051
rect 269869 20023 279237 20051
rect 279265 20023 279299 20051
rect 279327 20023 279361 20051
rect 279389 20023 279423 20051
rect 279451 20023 294597 20051
rect 294625 20023 294659 20051
rect 294687 20023 294721 20051
rect 294749 20023 294783 20051
rect 294811 20023 298248 20051
rect 298276 20023 298310 20051
rect 298338 20023 298372 20051
rect 298400 20023 298434 20051
rect 298462 20023 298990 20051
rect -958 19989 298990 20023
rect -958 19961 -430 19989
rect -402 19961 -368 19989
rect -340 19961 -306 19989
rect -278 19961 -244 19989
rect -216 19961 2757 19989
rect 2785 19961 2819 19989
rect 2847 19961 2881 19989
rect 2909 19961 2943 19989
rect 2971 19961 18117 19989
rect 18145 19961 18179 19989
rect 18207 19961 18241 19989
rect 18269 19961 18303 19989
rect 18331 19961 33477 19989
rect 33505 19961 33539 19989
rect 33567 19961 33601 19989
rect 33629 19961 33663 19989
rect 33691 19961 48837 19989
rect 48865 19961 48899 19989
rect 48927 19961 48961 19989
rect 48989 19961 49023 19989
rect 49051 19961 64197 19989
rect 64225 19961 64259 19989
rect 64287 19961 64321 19989
rect 64349 19961 64383 19989
rect 64411 19961 79557 19989
rect 79585 19961 79619 19989
rect 79647 19961 79681 19989
rect 79709 19961 79743 19989
rect 79771 19961 94917 19989
rect 94945 19961 94979 19989
rect 95007 19961 95041 19989
rect 95069 19961 95103 19989
rect 95131 19961 110277 19989
rect 110305 19961 110339 19989
rect 110367 19961 110401 19989
rect 110429 19961 110463 19989
rect 110491 19961 125637 19989
rect 125665 19961 125699 19989
rect 125727 19961 125761 19989
rect 125789 19961 125823 19989
rect 125851 19961 140997 19989
rect 141025 19961 141059 19989
rect 141087 19961 141121 19989
rect 141149 19961 141183 19989
rect 141211 19961 156357 19989
rect 156385 19961 156419 19989
rect 156447 19961 156481 19989
rect 156509 19961 156543 19989
rect 156571 19961 162259 19989
rect 162287 19961 162321 19989
rect 162349 19961 177619 19989
rect 177647 19961 177681 19989
rect 177709 19961 192979 19989
rect 193007 19961 193041 19989
rect 193069 19961 208339 19989
rect 208367 19961 208401 19989
rect 208429 19961 223699 19989
rect 223727 19961 223761 19989
rect 223789 19961 239059 19989
rect 239087 19961 239121 19989
rect 239149 19961 254419 19989
rect 254447 19961 254481 19989
rect 254509 19961 269779 19989
rect 269807 19961 269841 19989
rect 269869 19961 279237 19989
rect 279265 19961 279299 19989
rect 279327 19961 279361 19989
rect 279389 19961 279423 19989
rect 279451 19961 294597 19989
rect 294625 19961 294659 19989
rect 294687 19961 294721 19989
rect 294749 19961 294783 19989
rect 294811 19961 298248 19989
rect 298276 19961 298310 19989
rect 298338 19961 298372 19989
rect 298400 19961 298434 19989
rect 298462 19961 298990 19989
rect -958 19913 298990 19961
rect -958 14175 298990 14223
rect -958 14147 -910 14175
rect -882 14147 -848 14175
rect -820 14147 -786 14175
rect -758 14147 -724 14175
rect -696 14147 4617 14175
rect 4645 14147 4679 14175
rect 4707 14147 4741 14175
rect 4769 14147 4803 14175
rect 4831 14147 19977 14175
rect 20005 14147 20039 14175
rect 20067 14147 20101 14175
rect 20129 14147 20163 14175
rect 20191 14147 35337 14175
rect 35365 14147 35399 14175
rect 35427 14147 35461 14175
rect 35489 14147 35523 14175
rect 35551 14147 50697 14175
rect 50725 14147 50759 14175
rect 50787 14147 50821 14175
rect 50849 14147 50883 14175
rect 50911 14147 66057 14175
rect 66085 14147 66119 14175
rect 66147 14147 66181 14175
rect 66209 14147 66243 14175
rect 66271 14147 81417 14175
rect 81445 14147 81479 14175
rect 81507 14147 81541 14175
rect 81569 14147 81603 14175
rect 81631 14147 96777 14175
rect 96805 14147 96839 14175
rect 96867 14147 96901 14175
rect 96929 14147 96963 14175
rect 96991 14147 112137 14175
rect 112165 14147 112199 14175
rect 112227 14147 112261 14175
rect 112289 14147 112323 14175
rect 112351 14147 127497 14175
rect 127525 14147 127559 14175
rect 127587 14147 127621 14175
rect 127649 14147 127683 14175
rect 127711 14147 142857 14175
rect 142885 14147 142919 14175
rect 142947 14147 142981 14175
rect 143009 14147 143043 14175
rect 143071 14147 158217 14175
rect 158245 14147 158279 14175
rect 158307 14147 158341 14175
rect 158369 14147 158403 14175
rect 158431 14147 169939 14175
rect 169967 14147 170001 14175
rect 170029 14147 185299 14175
rect 185327 14147 185361 14175
rect 185389 14147 200659 14175
rect 200687 14147 200721 14175
rect 200749 14147 216019 14175
rect 216047 14147 216081 14175
rect 216109 14147 231379 14175
rect 231407 14147 231441 14175
rect 231469 14147 246739 14175
rect 246767 14147 246801 14175
rect 246829 14147 262099 14175
rect 262127 14147 262161 14175
rect 262189 14147 281097 14175
rect 281125 14147 281159 14175
rect 281187 14147 281221 14175
rect 281249 14147 281283 14175
rect 281311 14147 296457 14175
rect 296485 14147 296519 14175
rect 296547 14147 296581 14175
rect 296609 14147 296643 14175
rect 296671 14147 298728 14175
rect 298756 14147 298790 14175
rect 298818 14147 298852 14175
rect 298880 14147 298914 14175
rect 298942 14147 298990 14175
rect -958 14113 298990 14147
rect -958 14085 -910 14113
rect -882 14085 -848 14113
rect -820 14085 -786 14113
rect -758 14085 -724 14113
rect -696 14085 4617 14113
rect 4645 14085 4679 14113
rect 4707 14085 4741 14113
rect 4769 14085 4803 14113
rect 4831 14085 19977 14113
rect 20005 14085 20039 14113
rect 20067 14085 20101 14113
rect 20129 14085 20163 14113
rect 20191 14085 35337 14113
rect 35365 14085 35399 14113
rect 35427 14085 35461 14113
rect 35489 14085 35523 14113
rect 35551 14085 50697 14113
rect 50725 14085 50759 14113
rect 50787 14085 50821 14113
rect 50849 14085 50883 14113
rect 50911 14085 66057 14113
rect 66085 14085 66119 14113
rect 66147 14085 66181 14113
rect 66209 14085 66243 14113
rect 66271 14085 81417 14113
rect 81445 14085 81479 14113
rect 81507 14085 81541 14113
rect 81569 14085 81603 14113
rect 81631 14085 96777 14113
rect 96805 14085 96839 14113
rect 96867 14085 96901 14113
rect 96929 14085 96963 14113
rect 96991 14085 112137 14113
rect 112165 14085 112199 14113
rect 112227 14085 112261 14113
rect 112289 14085 112323 14113
rect 112351 14085 127497 14113
rect 127525 14085 127559 14113
rect 127587 14085 127621 14113
rect 127649 14085 127683 14113
rect 127711 14085 142857 14113
rect 142885 14085 142919 14113
rect 142947 14085 142981 14113
rect 143009 14085 143043 14113
rect 143071 14085 158217 14113
rect 158245 14085 158279 14113
rect 158307 14085 158341 14113
rect 158369 14085 158403 14113
rect 158431 14085 169939 14113
rect 169967 14085 170001 14113
rect 170029 14085 185299 14113
rect 185327 14085 185361 14113
rect 185389 14085 200659 14113
rect 200687 14085 200721 14113
rect 200749 14085 216019 14113
rect 216047 14085 216081 14113
rect 216109 14085 231379 14113
rect 231407 14085 231441 14113
rect 231469 14085 246739 14113
rect 246767 14085 246801 14113
rect 246829 14085 262099 14113
rect 262127 14085 262161 14113
rect 262189 14085 281097 14113
rect 281125 14085 281159 14113
rect 281187 14085 281221 14113
rect 281249 14085 281283 14113
rect 281311 14085 296457 14113
rect 296485 14085 296519 14113
rect 296547 14085 296581 14113
rect 296609 14085 296643 14113
rect 296671 14085 298728 14113
rect 298756 14085 298790 14113
rect 298818 14085 298852 14113
rect 298880 14085 298914 14113
rect 298942 14085 298990 14113
rect -958 14051 298990 14085
rect -958 14023 -910 14051
rect -882 14023 -848 14051
rect -820 14023 -786 14051
rect -758 14023 -724 14051
rect -696 14023 4617 14051
rect 4645 14023 4679 14051
rect 4707 14023 4741 14051
rect 4769 14023 4803 14051
rect 4831 14023 19977 14051
rect 20005 14023 20039 14051
rect 20067 14023 20101 14051
rect 20129 14023 20163 14051
rect 20191 14023 35337 14051
rect 35365 14023 35399 14051
rect 35427 14023 35461 14051
rect 35489 14023 35523 14051
rect 35551 14023 50697 14051
rect 50725 14023 50759 14051
rect 50787 14023 50821 14051
rect 50849 14023 50883 14051
rect 50911 14023 66057 14051
rect 66085 14023 66119 14051
rect 66147 14023 66181 14051
rect 66209 14023 66243 14051
rect 66271 14023 81417 14051
rect 81445 14023 81479 14051
rect 81507 14023 81541 14051
rect 81569 14023 81603 14051
rect 81631 14023 96777 14051
rect 96805 14023 96839 14051
rect 96867 14023 96901 14051
rect 96929 14023 96963 14051
rect 96991 14023 112137 14051
rect 112165 14023 112199 14051
rect 112227 14023 112261 14051
rect 112289 14023 112323 14051
rect 112351 14023 127497 14051
rect 127525 14023 127559 14051
rect 127587 14023 127621 14051
rect 127649 14023 127683 14051
rect 127711 14023 142857 14051
rect 142885 14023 142919 14051
rect 142947 14023 142981 14051
rect 143009 14023 143043 14051
rect 143071 14023 158217 14051
rect 158245 14023 158279 14051
rect 158307 14023 158341 14051
rect 158369 14023 158403 14051
rect 158431 14023 169939 14051
rect 169967 14023 170001 14051
rect 170029 14023 185299 14051
rect 185327 14023 185361 14051
rect 185389 14023 200659 14051
rect 200687 14023 200721 14051
rect 200749 14023 216019 14051
rect 216047 14023 216081 14051
rect 216109 14023 231379 14051
rect 231407 14023 231441 14051
rect 231469 14023 246739 14051
rect 246767 14023 246801 14051
rect 246829 14023 262099 14051
rect 262127 14023 262161 14051
rect 262189 14023 281097 14051
rect 281125 14023 281159 14051
rect 281187 14023 281221 14051
rect 281249 14023 281283 14051
rect 281311 14023 296457 14051
rect 296485 14023 296519 14051
rect 296547 14023 296581 14051
rect 296609 14023 296643 14051
rect 296671 14023 298728 14051
rect 298756 14023 298790 14051
rect 298818 14023 298852 14051
rect 298880 14023 298914 14051
rect 298942 14023 298990 14051
rect -958 13989 298990 14023
rect -958 13961 -910 13989
rect -882 13961 -848 13989
rect -820 13961 -786 13989
rect -758 13961 -724 13989
rect -696 13961 4617 13989
rect 4645 13961 4679 13989
rect 4707 13961 4741 13989
rect 4769 13961 4803 13989
rect 4831 13961 19977 13989
rect 20005 13961 20039 13989
rect 20067 13961 20101 13989
rect 20129 13961 20163 13989
rect 20191 13961 35337 13989
rect 35365 13961 35399 13989
rect 35427 13961 35461 13989
rect 35489 13961 35523 13989
rect 35551 13961 50697 13989
rect 50725 13961 50759 13989
rect 50787 13961 50821 13989
rect 50849 13961 50883 13989
rect 50911 13961 66057 13989
rect 66085 13961 66119 13989
rect 66147 13961 66181 13989
rect 66209 13961 66243 13989
rect 66271 13961 81417 13989
rect 81445 13961 81479 13989
rect 81507 13961 81541 13989
rect 81569 13961 81603 13989
rect 81631 13961 96777 13989
rect 96805 13961 96839 13989
rect 96867 13961 96901 13989
rect 96929 13961 96963 13989
rect 96991 13961 112137 13989
rect 112165 13961 112199 13989
rect 112227 13961 112261 13989
rect 112289 13961 112323 13989
rect 112351 13961 127497 13989
rect 127525 13961 127559 13989
rect 127587 13961 127621 13989
rect 127649 13961 127683 13989
rect 127711 13961 142857 13989
rect 142885 13961 142919 13989
rect 142947 13961 142981 13989
rect 143009 13961 143043 13989
rect 143071 13961 158217 13989
rect 158245 13961 158279 13989
rect 158307 13961 158341 13989
rect 158369 13961 158403 13989
rect 158431 13961 169939 13989
rect 169967 13961 170001 13989
rect 170029 13961 185299 13989
rect 185327 13961 185361 13989
rect 185389 13961 200659 13989
rect 200687 13961 200721 13989
rect 200749 13961 216019 13989
rect 216047 13961 216081 13989
rect 216109 13961 231379 13989
rect 231407 13961 231441 13989
rect 231469 13961 246739 13989
rect 246767 13961 246801 13989
rect 246829 13961 262099 13989
rect 262127 13961 262161 13989
rect 262189 13961 281097 13989
rect 281125 13961 281159 13989
rect 281187 13961 281221 13989
rect 281249 13961 281283 13989
rect 281311 13961 296457 13989
rect 296485 13961 296519 13989
rect 296547 13961 296581 13989
rect 296609 13961 296643 13989
rect 296671 13961 298728 13989
rect 298756 13961 298790 13989
rect 298818 13961 298852 13989
rect 298880 13961 298914 13989
rect 298942 13961 298990 13989
rect -958 13913 298990 13961
rect -958 11175 298990 11223
rect -958 11147 -430 11175
rect -402 11147 -368 11175
rect -340 11147 -306 11175
rect -278 11147 -244 11175
rect -216 11147 2757 11175
rect 2785 11147 2819 11175
rect 2847 11147 2881 11175
rect 2909 11147 2943 11175
rect 2971 11147 18117 11175
rect 18145 11147 18179 11175
rect 18207 11147 18241 11175
rect 18269 11147 18303 11175
rect 18331 11147 33477 11175
rect 33505 11147 33539 11175
rect 33567 11147 33601 11175
rect 33629 11147 33663 11175
rect 33691 11147 48837 11175
rect 48865 11147 48899 11175
rect 48927 11147 48961 11175
rect 48989 11147 49023 11175
rect 49051 11147 64197 11175
rect 64225 11147 64259 11175
rect 64287 11147 64321 11175
rect 64349 11147 64383 11175
rect 64411 11147 79557 11175
rect 79585 11147 79619 11175
rect 79647 11147 79681 11175
rect 79709 11147 79743 11175
rect 79771 11147 94917 11175
rect 94945 11147 94979 11175
rect 95007 11147 95041 11175
rect 95069 11147 95103 11175
rect 95131 11147 110277 11175
rect 110305 11147 110339 11175
rect 110367 11147 110401 11175
rect 110429 11147 110463 11175
rect 110491 11147 125637 11175
rect 125665 11147 125699 11175
rect 125727 11147 125761 11175
rect 125789 11147 125823 11175
rect 125851 11147 140997 11175
rect 141025 11147 141059 11175
rect 141087 11147 141121 11175
rect 141149 11147 141183 11175
rect 141211 11147 156357 11175
rect 156385 11147 156419 11175
rect 156447 11147 156481 11175
rect 156509 11147 156543 11175
rect 156571 11147 162259 11175
rect 162287 11147 162321 11175
rect 162349 11147 177619 11175
rect 177647 11147 177681 11175
rect 177709 11147 192979 11175
rect 193007 11147 193041 11175
rect 193069 11147 208339 11175
rect 208367 11147 208401 11175
rect 208429 11147 223699 11175
rect 223727 11147 223761 11175
rect 223789 11147 239059 11175
rect 239087 11147 239121 11175
rect 239149 11147 254419 11175
rect 254447 11147 254481 11175
rect 254509 11147 269779 11175
rect 269807 11147 269841 11175
rect 269869 11147 279237 11175
rect 279265 11147 279299 11175
rect 279327 11147 279361 11175
rect 279389 11147 279423 11175
rect 279451 11147 294597 11175
rect 294625 11147 294659 11175
rect 294687 11147 294721 11175
rect 294749 11147 294783 11175
rect 294811 11147 298248 11175
rect 298276 11147 298310 11175
rect 298338 11147 298372 11175
rect 298400 11147 298434 11175
rect 298462 11147 298990 11175
rect -958 11113 298990 11147
rect -958 11085 -430 11113
rect -402 11085 -368 11113
rect -340 11085 -306 11113
rect -278 11085 -244 11113
rect -216 11085 2757 11113
rect 2785 11085 2819 11113
rect 2847 11085 2881 11113
rect 2909 11085 2943 11113
rect 2971 11085 18117 11113
rect 18145 11085 18179 11113
rect 18207 11085 18241 11113
rect 18269 11085 18303 11113
rect 18331 11085 33477 11113
rect 33505 11085 33539 11113
rect 33567 11085 33601 11113
rect 33629 11085 33663 11113
rect 33691 11085 48837 11113
rect 48865 11085 48899 11113
rect 48927 11085 48961 11113
rect 48989 11085 49023 11113
rect 49051 11085 64197 11113
rect 64225 11085 64259 11113
rect 64287 11085 64321 11113
rect 64349 11085 64383 11113
rect 64411 11085 79557 11113
rect 79585 11085 79619 11113
rect 79647 11085 79681 11113
rect 79709 11085 79743 11113
rect 79771 11085 94917 11113
rect 94945 11085 94979 11113
rect 95007 11085 95041 11113
rect 95069 11085 95103 11113
rect 95131 11085 110277 11113
rect 110305 11085 110339 11113
rect 110367 11085 110401 11113
rect 110429 11085 110463 11113
rect 110491 11085 125637 11113
rect 125665 11085 125699 11113
rect 125727 11085 125761 11113
rect 125789 11085 125823 11113
rect 125851 11085 140997 11113
rect 141025 11085 141059 11113
rect 141087 11085 141121 11113
rect 141149 11085 141183 11113
rect 141211 11085 156357 11113
rect 156385 11085 156419 11113
rect 156447 11085 156481 11113
rect 156509 11085 156543 11113
rect 156571 11085 162259 11113
rect 162287 11085 162321 11113
rect 162349 11085 177619 11113
rect 177647 11085 177681 11113
rect 177709 11085 192979 11113
rect 193007 11085 193041 11113
rect 193069 11085 208339 11113
rect 208367 11085 208401 11113
rect 208429 11085 223699 11113
rect 223727 11085 223761 11113
rect 223789 11085 239059 11113
rect 239087 11085 239121 11113
rect 239149 11085 254419 11113
rect 254447 11085 254481 11113
rect 254509 11085 269779 11113
rect 269807 11085 269841 11113
rect 269869 11085 279237 11113
rect 279265 11085 279299 11113
rect 279327 11085 279361 11113
rect 279389 11085 279423 11113
rect 279451 11085 294597 11113
rect 294625 11085 294659 11113
rect 294687 11085 294721 11113
rect 294749 11085 294783 11113
rect 294811 11085 298248 11113
rect 298276 11085 298310 11113
rect 298338 11085 298372 11113
rect 298400 11085 298434 11113
rect 298462 11085 298990 11113
rect -958 11051 298990 11085
rect -958 11023 -430 11051
rect -402 11023 -368 11051
rect -340 11023 -306 11051
rect -278 11023 -244 11051
rect -216 11023 2757 11051
rect 2785 11023 2819 11051
rect 2847 11023 2881 11051
rect 2909 11023 2943 11051
rect 2971 11023 18117 11051
rect 18145 11023 18179 11051
rect 18207 11023 18241 11051
rect 18269 11023 18303 11051
rect 18331 11023 33477 11051
rect 33505 11023 33539 11051
rect 33567 11023 33601 11051
rect 33629 11023 33663 11051
rect 33691 11023 48837 11051
rect 48865 11023 48899 11051
rect 48927 11023 48961 11051
rect 48989 11023 49023 11051
rect 49051 11023 64197 11051
rect 64225 11023 64259 11051
rect 64287 11023 64321 11051
rect 64349 11023 64383 11051
rect 64411 11023 79557 11051
rect 79585 11023 79619 11051
rect 79647 11023 79681 11051
rect 79709 11023 79743 11051
rect 79771 11023 94917 11051
rect 94945 11023 94979 11051
rect 95007 11023 95041 11051
rect 95069 11023 95103 11051
rect 95131 11023 110277 11051
rect 110305 11023 110339 11051
rect 110367 11023 110401 11051
rect 110429 11023 110463 11051
rect 110491 11023 125637 11051
rect 125665 11023 125699 11051
rect 125727 11023 125761 11051
rect 125789 11023 125823 11051
rect 125851 11023 140997 11051
rect 141025 11023 141059 11051
rect 141087 11023 141121 11051
rect 141149 11023 141183 11051
rect 141211 11023 156357 11051
rect 156385 11023 156419 11051
rect 156447 11023 156481 11051
rect 156509 11023 156543 11051
rect 156571 11023 162259 11051
rect 162287 11023 162321 11051
rect 162349 11023 177619 11051
rect 177647 11023 177681 11051
rect 177709 11023 192979 11051
rect 193007 11023 193041 11051
rect 193069 11023 208339 11051
rect 208367 11023 208401 11051
rect 208429 11023 223699 11051
rect 223727 11023 223761 11051
rect 223789 11023 239059 11051
rect 239087 11023 239121 11051
rect 239149 11023 254419 11051
rect 254447 11023 254481 11051
rect 254509 11023 269779 11051
rect 269807 11023 269841 11051
rect 269869 11023 279237 11051
rect 279265 11023 279299 11051
rect 279327 11023 279361 11051
rect 279389 11023 279423 11051
rect 279451 11023 294597 11051
rect 294625 11023 294659 11051
rect 294687 11023 294721 11051
rect 294749 11023 294783 11051
rect 294811 11023 298248 11051
rect 298276 11023 298310 11051
rect 298338 11023 298372 11051
rect 298400 11023 298434 11051
rect 298462 11023 298990 11051
rect -958 10989 298990 11023
rect -958 10961 -430 10989
rect -402 10961 -368 10989
rect -340 10961 -306 10989
rect -278 10961 -244 10989
rect -216 10961 2757 10989
rect 2785 10961 2819 10989
rect 2847 10961 2881 10989
rect 2909 10961 2943 10989
rect 2971 10961 18117 10989
rect 18145 10961 18179 10989
rect 18207 10961 18241 10989
rect 18269 10961 18303 10989
rect 18331 10961 33477 10989
rect 33505 10961 33539 10989
rect 33567 10961 33601 10989
rect 33629 10961 33663 10989
rect 33691 10961 48837 10989
rect 48865 10961 48899 10989
rect 48927 10961 48961 10989
rect 48989 10961 49023 10989
rect 49051 10961 64197 10989
rect 64225 10961 64259 10989
rect 64287 10961 64321 10989
rect 64349 10961 64383 10989
rect 64411 10961 79557 10989
rect 79585 10961 79619 10989
rect 79647 10961 79681 10989
rect 79709 10961 79743 10989
rect 79771 10961 94917 10989
rect 94945 10961 94979 10989
rect 95007 10961 95041 10989
rect 95069 10961 95103 10989
rect 95131 10961 110277 10989
rect 110305 10961 110339 10989
rect 110367 10961 110401 10989
rect 110429 10961 110463 10989
rect 110491 10961 125637 10989
rect 125665 10961 125699 10989
rect 125727 10961 125761 10989
rect 125789 10961 125823 10989
rect 125851 10961 140997 10989
rect 141025 10961 141059 10989
rect 141087 10961 141121 10989
rect 141149 10961 141183 10989
rect 141211 10961 156357 10989
rect 156385 10961 156419 10989
rect 156447 10961 156481 10989
rect 156509 10961 156543 10989
rect 156571 10961 162259 10989
rect 162287 10961 162321 10989
rect 162349 10961 177619 10989
rect 177647 10961 177681 10989
rect 177709 10961 192979 10989
rect 193007 10961 193041 10989
rect 193069 10961 208339 10989
rect 208367 10961 208401 10989
rect 208429 10961 223699 10989
rect 223727 10961 223761 10989
rect 223789 10961 239059 10989
rect 239087 10961 239121 10989
rect 239149 10961 254419 10989
rect 254447 10961 254481 10989
rect 254509 10961 269779 10989
rect 269807 10961 269841 10989
rect 269869 10961 279237 10989
rect 279265 10961 279299 10989
rect 279327 10961 279361 10989
rect 279389 10961 279423 10989
rect 279451 10961 294597 10989
rect 294625 10961 294659 10989
rect 294687 10961 294721 10989
rect 294749 10961 294783 10989
rect 294811 10961 298248 10989
rect 298276 10961 298310 10989
rect 298338 10961 298372 10989
rect 298400 10961 298434 10989
rect 298462 10961 298990 10989
rect -958 10913 298990 10961
rect -958 5175 298990 5223
rect -958 5147 -910 5175
rect -882 5147 -848 5175
rect -820 5147 -786 5175
rect -758 5147 -724 5175
rect -696 5147 4617 5175
rect 4645 5147 4679 5175
rect 4707 5147 4741 5175
rect 4769 5147 4803 5175
rect 4831 5147 19977 5175
rect 20005 5147 20039 5175
rect 20067 5147 20101 5175
rect 20129 5147 20163 5175
rect 20191 5147 35337 5175
rect 35365 5147 35399 5175
rect 35427 5147 35461 5175
rect 35489 5147 35523 5175
rect 35551 5147 50697 5175
rect 50725 5147 50759 5175
rect 50787 5147 50821 5175
rect 50849 5147 50883 5175
rect 50911 5147 66057 5175
rect 66085 5147 66119 5175
rect 66147 5147 66181 5175
rect 66209 5147 66243 5175
rect 66271 5147 81417 5175
rect 81445 5147 81479 5175
rect 81507 5147 81541 5175
rect 81569 5147 81603 5175
rect 81631 5147 96777 5175
rect 96805 5147 96839 5175
rect 96867 5147 96901 5175
rect 96929 5147 96963 5175
rect 96991 5147 112137 5175
rect 112165 5147 112199 5175
rect 112227 5147 112261 5175
rect 112289 5147 112323 5175
rect 112351 5147 127497 5175
rect 127525 5147 127559 5175
rect 127587 5147 127621 5175
rect 127649 5147 127683 5175
rect 127711 5147 142857 5175
rect 142885 5147 142919 5175
rect 142947 5147 142981 5175
rect 143009 5147 143043 5175
rect 143071 5147 158217 5175
rect 158245 5147 158279 5175
rect 158307 5147 158341 5175
rect 158369 5147 158403 5175
rect 158431 5147 173577 5175
rect 173605 5147 173639 5175
rect 173667 5147 173701 5175
rect 173729 5147 173763 5175
rect 173791 5147 188937 5175
rect 188965 5147 188999 5175
rect 189027 5147 189061 5175
rect 189089 5147 189123 5175
rect 189151 5147 204297 5175
rect 204325 5147 204359 5175
rect 204387 5147 204421 5175
rect 204449 5147 204483 5175
rect 204511 5147 219657 5175
rect 219685 5147 219719 5175
rect 219747 5147 219781 5175
rect 219809 5147 219843 5175
rect 219871 5147 235017 5175
rect 235045 5147 235079 5175
rect 235107 5147 235141 5175
rect 235169 5147 235203 5175
rect 235231 5147 250377 5175
rect 250405 5147 250439 5175
rect 250467 5147 250501 5175
rect 250529 5147 250563 5175
rect 250591 5147 265737 5175
rect 265765 5147 265799 5175
rect 265827 5147 265861 5175
rect 265889 5147 265923 5175
rect 265951 5147 281097 5175
rect 281125 5147 281159 5175
rect 281187 5147 281221 5175
rect 281249 5147 281283 5175
rect 281311 5147 296457 5175
rect 296485 5147 296519 5175
rect 296547 5147 296581 5175
rect 296609 5147 296643 5175
rect 296671 5147 298728 5175
rect 298756 5147 298790 5175
rect 298818 5147 298852 5175
rect 298880 5147 298914 5175
rect 298942 5147 298990 5175
rect -958 5113 298990 5147
rect -958 5085 -910 5113
rect -882 5085 -848 5113
rect -820 5085 -786 5113
rect -758 5085 -724 5113
rect -696 5085 4617 5113
rect 4645 5085 4679 5113
rect 4707 5085 4741 5113
rect 4769 5085 4803 5113
rect 4831 5085 19977 5113
rect 20005 5085 20039 5113
rect 20067 5085 20101 5113
rect 20129 5085 20163 5113
rect 20191 5085 35337 5113
rect 35365 5085 35399 5113
rect 35427 5085 35461 5113
rect 35489 5085 35523 5113
rect 35551 5085 50697 5113
rect 50725 5085 50759 5113
rect 50787 5085 50821 5113
rect 50849 5085 50883 5113
rect 50911 5085 66057 5113
rect 66085 5085 66119 5113
rect 66147 5085 66181 5113
rect 66209 5085 66243 5113
rect 66271 5085 81417 5113
rect 81445 5085 81479 5113
rect 81507 5085 81541 5113
rect 81569 5085 81603 5113
rect 81631 5085 96777 5113
rect 96805 5085 96839 5113
rect 96867 5085 96901 5113
rect 96929 5085 96963 5113
rect 96991 5085 112137 5113
rect 112165 5085 112199 5113
rect 112227 5085 112261 5113
rect 112289 5085 112323 5113
rect 112351 5085 127497 5113
rect 127525 5085 127559 5113
rect 127587 5085 127621 5113
rect 127649 5085 127683 5113
rect 127711 5085 142857 5113
rect 142885 5085 142919 5113
rect 142947 5085 142981 5113
rect 143009 5085 143043 5113
rect 143071 5085 158217 5113
rect 158245 5085 158279 5113
rect 158307 5085 158341 5113
rect 158369 5085 158403 5113
rect 158431 5085 173577 5113
rect 173605 5085 173639 5113
rect 173667 5085 173701 5113
rect 173729 5085 173763 5113
rect 173791 5085 188937 5113
rect 188965 5085 188999 5113
rect 189027 5085 189061 5113
rect 189089 5085 189123 5113
rect 189151 5085 204297 5113
rect 204325 5085 204359 5113
rect 204387 5085 204421 5113
rect 204449 5085 204483 5113
rect 204511 5085 219657 5113
rect 219685 5085 219719 5113
rect 219747 5085 219781 5113
rect 219809 5085 219843 5113
rect 219871 5085 235017 5113
rect 235045 5085 235079 5113
rect 235107 5085 235141 5113
rect 235169 5085 235203 5113
rect 235231 5085 250377 5113
rect 250405 5085 250439 5113
rect 250467 5085 250501 5113
rect 250529 5085 250563 5113
rect 250591 5085 265737 5113
rect 265765 5085 265799 5113
rect 265827 5085 265861 5113
rect 265889 5085 265923 5113
rect 265951 5085 281097 5113
rect 281125 5085 281159 5113
rect 281187 5085 281221 5113
rect 281249 5085 281283 5113
rect 281311 5085 296457 5113
rect 296485 5085 296519 5113
rect 296547 5085 296581 5113
rect 296609 5085 296643 5113
rect 296671 5085 298728 5113
rect 298756 5085 298790 5113
rect 298818 5085 298852 5113
rect 298880 5085 298914 5113
rect 298942 5085 298990 5113
rect -958 5051 298990 5085
rect -958 5023 -910 5051
rect -882 5023 -848 5051
rect -820 5023 -786 5051
rect -758 5023 -724 5051
rect -696 5023 4617 5051
rect 4645 5023 4679 5051
rect 4707 5023 4741 5051
rect 4769 5023 4803 5051
rect 4831 5023 19977 5051
rect 20005 5023 20039 5051
rect 20067 5023 20101 5051
rect 20129 5023 20163 5051
rect 20191 5023 35337 5051
rect 35365 5023 35399 5051
rect 35427 5023 35461 5051
rect 35489 5023 35523 5051
rect 35551 5023 50697 5051
rect 50725 5023 50759 5051
rect 50787 5023 50821 5051
rect 50849 5023 50883 5051
rect 50911 5023 66057 5051
rect 66085 5023 66119 5051
rect 66147 5023 66181 5051
rect 66209 5023 66243 5051
rect 66271 5023 81417 5051
rect 81445 5023 81479 5051
rect 81507 5023 81541 5051
rect 81569 5023 81603 5051
rect 81631 5023 96777 5051
rect 96805 5023 96839 5051
rect 96867 5023 96901 5051
rect 96929 5023 96963 5051
rect 96991 5023 112137 5051
rect 112165 5023 112199 5051
rect 112227 5023 112261 5051
rect 112289 5023 112323 5051
rect 112351 5023 127497 5051
rect 127525 5023 127559 5051
rect 127587 5023 127621 5051
rect 127649 5023 127683 5051
rect 127711 5023 142857 5051
rect 142885 5023 142919 5051
rect 142947 5023 142981 5051
rect 143009 5023 143043 5051
rect 143071 5023 158217 5051
rect 158245 5023 158279 5051
rect 158307 5023 158341 5051
rect 158369 5023 158403 5051
rect 158431 5023 173577 5051
rect 173605 5023 173639 5051
rect 173667 5023 173701 5051
rect 173729 5023 173763 5051
rect 173791 5023 188937 5051
rect 188965 5023 188999 5051
rect 189027 5023 189061 5051
rect 189089 5023 189123 5051
rect 189151 5023 204297 5051
rect 204325 5023 204359 5051
rect 204387 5023 204421 5051
rect 204449 5023 204483 5051
rect 204511 5023 219657 5051
rect 219685 5023 219719 5051
rect 219747 5023 219781 5051
rect 219809 5023 219843 5051
rect 219871 5023 235017 5051
rect 235045 5023 235079 5051
rect 235107 5023 235141 5051
rect 235169 5023 235203 5051
rect 235231 5023 250377 5051
rect 250405 5023 250439 5051
rect 250467 5023 250501 5051
rect 250529 5023 250563 5051
rect 250591 5023 265737 5051
rect 265765 5023 265799 5051
rect 265827 5023 265861 5051
rect 265889 5023 265923 5051
rect 265951 5023 281097 5051
rect 281125 5023 281159 5051
rect 281187 5023 281221 5051
rect 281249 5023 281283 5051
rect 281311 5023 296457 5051
rect 296485 5023 296519 5051
rect 296547 5023 296581 5051
rect 296609 5023 296643 5051
rect 296671 5023 298728 5051
rect 298756 5023 298790 5051
rect 298818 5023 298852 5051
rect 298880 5023 298914 5051
rect 298942 5023 298990 5051
rect -958 4989 298990 5023
rect -958 4961 -910 4989
rect -882 4961 -848 4989
rect -820 4961 -786 4989
rect -758 4961 -724 4989
rect -696 4961 4617 4989
rect 4645 4961 4679 4989
rect 4707 4961 4741 4989
rect 4769 4961 4803 4989
rect 4831 4961 19977 4989
rect 20005 4961 20039 4989
rect 20067 4961 20101 4989
rect 20129 4961 20163 4989
rect 20191 4961 35337 4989
rect 35365 4961 35399 4989
rect 35427 4961 35461 4989
rect 35489 4961 35523 4989
rect 35551 4961 50697 4989
rect 50725 4961 50759 4989
rect 50787 4961 50821 4989
rect 50849 4961 50883 4989
rect 50911 4961 66057 4989
rect 66085 4961 66119 4989
rect 66147 4961 66181 4989
rect 66209 4961 66243 4989
rect 66271 4961 81417 4989
rect 81445 4961 81479 4989
rect 81507 4961 81541 4989
rect 81569 4961 81603 4989
rect 81631 4961 96777 4989
rect 96805 4961 96839 4989
rect 96867 4961 96901 4989
rect 96929 4961 96963 4989
rect 96991 4961 112137 4989
rect 112165 4961 112199 4989
rect 112227 4961 112261 4989
rect 112289 4961 112323 4989
rect 112351 4961 127497 4989
rect 127525 4961 127559 4989
rect 127587 4961 127621 4989
rect 127649 4961 127683 4989
rect 127711 4961 142857 4989
rect 142885 4961 142919 4989
rect 142947 4961 142981 4989
rect 143009 4961 143043 4989
rect 143071 4961 158217 4989
rect 158245 4961 158279 4989
rect 158307 4961 158341 4989
rect 158369 4961 158403 4989
rect 158431 4961 173577 4989
rect 173605 4961 173639 4989
rect 173667 4961 173701 4989
rect 173729 4961 173763 4989
rect 173791 4961 188937 4989
rect 188965 4961 188999 4989
rect 189027 4961 189061 4989
rect 189089 4961 189123 4989
rect 189151 4961 204297 4989
rect 204325 4961 204359 4989
rect 204387 4961 204421 4989
rect 204449 4961 204483 4989
rect 204511 4961 219657 4989
rect 219685 4961 219719 4989
rect 219747 4961 219781 4989
rect 219809 4961 219843 4989
rect 219871 4961 235017 4989
rect 235045 4961 235079 4989
rect 235107 4961 235141 4989
rect 235169 4961 235203 4989
rect 235231 4961 250377 4989
rect 250405 4961 250439 4989
rect 250467 4961 250501 4989
rect 250529 4961 250563 4989
rect 250591 4961 265737 4989
rect 265765 4961 265799 4989
rect 265827 4961 265861 4989
rect 265889 4961 265923 4989
rect 265951 4961 281097 4989
rect 281125 4961 281159 4989
rect 281187 4961 281221 4989
rect 281249 4961 281283 4989
rect 281311 4961 296457 4989
rect 296485 4961 296519 4989
rect 296547 4961 296581 4989
rect 296609 4961 296643 4989
rect 296671 4961 298728 4989
rect 298756 4961 298790 4989
rect 298818 4961 298852 4989
rect 298880 4961 298914 4989
rect 298942 4961 298990 4989
rect -958 4913 298990 4961
rect -958 2175 298990 2223
rect -958 2147 -430 2175
rect -402 2147 -368 2175
rect -340 2147 -306 2175
rect -278 2147 -244 2175
rect -216 2147 2757 2175
rect 2785 2147 2819 2175
rect 2847 2147 2881 2175
rect 2909 2147 2943 2175
rect 2971 2147 18117 2175
rect 18145 2147 18179 2175
rect 18207 2147 18241 2175
rect 18269 2147 18303 2175
rect 18331 2147 33477 2175
rect 33505 2147 33539 2175
rect 33567 2147 33601 2175
rect 33629 2147 33663 2175
rect 33691 2147 48837 2175
rect 48865 2147 48899 2175
rect 48927 2147 48961 2175
rect 48989 2147 49023 2175
rect 49051 2147 64197 2175
rect 64225 2147 64259 2175
rect 64287 2147 64321 2175
rect 64349 2147 64383 2175
rect 64411 2147 79557 2175
rect 79585 2147 79619 2175
rect 79647 2147 79681 2175
rect 79709 2147 79743 2175
rect 79771 2147 94917 2175
rect 94945 2147 94979 2175
rect 95007 2147 95041 2175
rect 95069 2147 95103 2175
rect 95131 2147 110277 2175
rect 110305 2147 110339 2175
rect 110367 2147 110401 2175
rect 110429 2147 110463 2175
rect 110491 2147 125637 2175
rect 125665 2147 125699 2175
rect 125727 2147 125761 2175
rect 125789 2147 125823 2175
rect 125851 2147 140997 2175
rect 141025 2147 141059 2175
rect 141087 2147 141121 2175
rect 141149 2147 141183 2175
rect 141211 2147 156357 2175
rect 156385 2147 156419 2175
rect 156447 2147 156481 2175
rect 156509 2147 156543 2175
rect 156571 2147 171717 2175
rect 171745 2147 171779 2175
rect 171807 2147 171841 2175
rect 171869 2147 171903 2175
rect 171931 2147 187077 2175
rect 187105 2147 187139 2175
rect 187167 2147 187201 2175
rect 187229 2147 187263 2175
rect 187291 2147 202437 2175
rect 202465 2147 202499 2175
rect 202527 2147 202561 2175
rect 202589 2147 202623 2175
rect 202651 2147 217797 2175
rect 217825 2147 217859 2175
rect 217887 2147 217921 2175
rect 217949 2147 217983 2175
rect 218011 2147 233157 2175
rect 233185 2147 233219 2175
rect 233247 2147 233281 2175
rect 233309 2147 233343 2175
rect 233371 2147 248517 2175
rect 248545 2147 248579 2175
rect 248607 2147 248641 2175
rect 248669 2147 248703 2175
rect 248731 2147 263877 2175
rect 263905 2147 263939 2175
rect 263967 2147 264001 2175
rect 264029 2147 264063 2175
rect 264091 2147 279237 2175
rect 279265 2147 279299 2175
rect 279327 2147 279361 2175
rect 279389 2147 279423 2175
rect 279451 2147 294597 2175
rect 294625 2147 294659 2175
rect 294687 2147 294721 2175
rect 294749 2147 294783 2175
rect 294811 2147 298248 2175
rect 298276 2147 298310 2175
rect 298338 2147 298372 2175
rect 298400 2147 298434 2175
rect 298462 2147 298990 2175
rect -958 2113 298990 2147
rect -958 2085 -430 2113
rect -402 2085 -368 2113
rect -340 2085 -306 2113
rect -278 2085 -244 2113
rect -216 2085 2757 2113
rect 2785 2085 2819 2113
rect 2847 2085 2881 2113
rect 2909 2085 2943 2113
rect 2971 2085 18117 2113
rect 18145 2085 18179 2113
rect 18207 2085 18241 2113
rect 18269 2085 18303 2113
rect 18331 2085 33477 2113
rect 33505 2085 33539 2113
rect 33567 2085 33601 2113
rect 33629 2085 33663 2113
rect 33691 2085 48837 2113
rect 48865 2085 48899 2113
rect 48927 2085 48961 2113
rect 48989 2085 49023 2113
rect 49051 2085 64197 2113
rect 64225 2085 64259 2113
rect 64287 2085 64321 2113
rect 64349 2085 64383 2113
rect 64411 2085 79557 2113
rect 79585 2085 79619 2113
rect 79647 2085 79681 2113
rect 79709 2085 79743 2113
rect 79771 2085 94917 2113
rect 94945 2085 94979 2113
rect 95007 2085 95041 2113
rect 95069 2085 95103 2113
rect 95131 2085 110277 2113
rect 110305 2085 110339 2113
rect 110367 2085 110401 2113
rect 110429 2085 110463 2113
rect 110491 2085 125637 2113
rect 125665 2085 125699 2113
rect 125727 2085 125761 2113
rect 125789 2085 125823 2113
rect 125851 2085 140997 2113
rect 141025 2085 141059 2113
rect 141087 2085 141121 2113
rect 141149 2085 141183 2113
rect 141211 2085 156357 2113
rect 156385 2085 156419 2113
rect 156447 2085 156481 2113
rect 156509 2085 156543 2113
rect 156571 2085 171717 2113
rect 171745 2085 171779 2113
rect 171807 2085 171841 2113
rect 171869 2085 171903 2113
rect 171931 2085 187077 2113
rect 187105 2085 187139 2113
rect 187167 2085 187201 2113
rect 187229 2085 187263 2113
rect 187291 2085 202437 2113
rect 202465 2085 202499 2113
rect 202527 2085 202561 2113
rect 202589 2085 202623 2113
rect 202651 2085 217797 2113
rect 217825 2085 217859 2113
rect 217887 2085 217921 2113
rect 217949 2085 217983 2113
rect 218011 2085 233157 2113
rect 233185 2085 233219 2113
rect 233247 2085 233281 2113
rect 233309 2085 233343 2113
rect 233371 2085 248517 2113
rect 248545 2085 248579 2113
rect 248607 2085 248641 2113
rect 248669 2085 248703 2113
rect 248731 2085 263877 2113
rect 263905 2085 263939 2113
rect 263967 2085 264001 2113
rect 264029 2085 264063 2113
rect 264091 2085 279237 2113
rect 279265 2085 279299 2113
rect 279327 2085 279361 2113
rect 279389 2085 279423 2113
rect 279451 2085 294597 2113
rect 294625 2085 294659 2113
rect 294687 2085 294721 2113
rect 294749 2085 294783 2113
rect 294811 2085 298248 2113
rect 298276 2085 298310 2113
rect 298338 2085 298372 2113
rect 298400 2085 298434 2113
rect 298462 2085 298990 2113
rect -958 2051 298990 2085
rect -958 2023 -430 2051
rect -402 2023 -368 2051
rect -340 2023 -306 2051
rect -278 2023 -244 2051
rect -216 2023 2757 2051
rect 2785 2023 2819 2051
rect 2847 2023 2881 2051
rect 2909 2023 2943 2051
rect 2971 2023 18117 2051
rect 18145 2023 18179 2051
rect 18207 2023 18241 2051
rect 18269 2023 18303 2051
rect 18331 2023 33477 2051
rect 33505 2023 33539 2051
rect 33567 2023 33601 2051
rect 33629 2023 33663 2051
rect 33691 2023 48837 2051
rect 48865 2023 48899 2051
rect 48927 2023 48961 2051
rect 48989 2023 49023 2051
rect 49051 2023 64197 2051
rect 64225 2023 64259 2051
rect 64287 2023 64321 2051
rect 64349 2023 64383 2051
rect 64411 2023 79557 2051
rect 79585 2023 79619 2051
rect 79647 2023 79681 2051
rect 79709 2023 79743 2051
rect 79771 2023 94917 2051
rect 94945 2023 94979 2051
rect 95007 2023 95041 2051
rect 95069 2023 95103 2051
rect 95131 2023 110277 2051
rect 110305 2023 110339 2051
rect 110367 2023 110401 2051
rect 110429 2023 110463 2051
rect 110491 2023 125637 2051
rect 125665 2023 125699 2051
rect 125727 2023 125761 2051
rect 125789 2023 125823 2051
rect 125851 2023 140997 2051
rect 141025 2023 141059 2051
rect 141087 2023 141121 2051
rect 141149 2023 141183 2051
rect 141211 2023 156357 2051
rect 156385 2023 156419 2051
rect 156447 2023 156481 2051
rect 156509 2023 156543 2051
rect 156571 2023 171717 2051
rect 171745 2023 171779 2051
rect 171807 2023 171841 2051
rect 171869 2023 171903 2051
rect 171931 2023 187077 2051
rect 187105 2023 187139 2051
rect 187167 2023 187201 2051
rect 187229 2023 187263 2051
rect 187291 2023 202437 2051
rect 202465 2023 202499 2051
rect 202527 2023 202561 2051
rect 202589 2023 202623 2051
rect 202651 2023 217797 2051
rect 217825 2023 217859 2051
rect 217887 2023 217921 2051
rect 217949 2023 217983 2051
rect 218011 2023 233157 2051
rect 233185 2023 233219 2051
rect 233247 2023 233281 2051
rect 233309 2023 233343 2051
rect 233371 2023 248517 2051
rect 248545 2023 248579 2051
rect 248607 2023 248641 2051
rect 248669 2023 248703 2051
rect 248731 2023 263877 2051
rect 263905 2023 263939 2051
rect 263967 2023 264001 2051
rect 264029 2023 264063 2051
rect 264091 2023 279237 2051
rect 279265 2023 279299 2051
rect 279327 2023 279361 2051
rect 279389 2023 279423 2051
rect 279451 2023 294597 2051
rect 294625 2023 294659 2051
rect 294687 2023 294721 2051
rect 294749 2023 294783 2051
rect 294811 2023 298248 2051
rect 298276 2023 298310 2051
rect 298338 2023 298372 2051
rect 298400 2023 298434 2051
rect 298462 2023 298990 2051
rect -958 1989 298990 2023
rect -958 1961 -430 1989
rect -402 1961 -368 1989
rect -340 1961 -306 1989
rect -278 1961 -244 1989
rect -216 1961 2757 1989
rect 2785 1961 2819 1989
rect 2847 1961 2881 1989
rect 2909 1961 2943 1989
rect 2971 1961 18117 1989
rect 18145 1961 18179 1989
rect 18207 1961 18241 1989
rect 18269 1961 18303 1989
rect 18331 1961 33477 1989
rect 33505 1961 33539 1989
rect 33567 1961 33601 1989
rect 33629 1961 33663 1989
rect 33691 1961 48837 1989
rect 48865 1961 48899 1989
rect 48927 1961 48961 1989
rect 48989 1961 49023 1989
rect 49051 1961 64197 1989
rect 64225 1961 64259 1989
rect 64287 1961 64321 1989
rect 64349 1961 64383 1989
rect 64411 1961 79557 1989
rect 79585 1961 79619 1989
rect 79647 1961 79681 1989
rect 79709 1961 79743 1989
rect 79771 1961 94917 1989
rect 94945 1961 94979 1989
rect 95007 1961 95041 1989
rect 95069 1961 95103 1989
rect 95131 1961 110277 1989
rect 110305 1961 110339 1989
rect 110367 1961 110401 1989
rect 110429 1961 110463 1989
rect 110491 1961 125637 1989
rect 125665 1961 125699 1989
rect 125727 1961 125761 1989
rect 125789 1961 125823 1989
rect 125851 1961 140997 1989
rect 141025 1961 141059 1989
rect 141087 1961 141121 1989
rect 141149 1961 141183 1989
rect 141211 1961 156357 1989
rect 156385 1961 156419 1989
rect 156447 1961 156481 1989
rect 156509 1961 156543 1989
rect 156571 1961 171717 1989
rect 171745 1961 171779 1989
rect 171807 1961 171841 1989
rect 171869 1961 171903 1989
rect 171931 1961 187077 1989
rect 187105 1961 187139 1989
rect 187167 1961 187201 1989
rect 187229 1961 187263 1989
rect 187291 1961 202437 1989
rect 202465 1961 202499 1989
rect 202527 1961 202561 1989
rect 202589 1961 202623 1989
rect 202651 1961 217797 1989
rect 217825 1961 217859 1989
rect 217887 1961 217921 1989
rect 217949 1961 217983 1989
rect 218011 1961 233157 1989
rect 233185 1961 233219 1989
rect 233247 1961 233281 1989
rect 233309 1961 233343 1989
rect 233371 1961 248517 1989
rect 248545 1961 248579 1989
rect 248607 1961 248641 1989
rect 248669 1961 248703 1989
rect 248731 1961 263877 1989
rect 263905 1961 263939 1989
rect 263967 1961 264001 1989
rect 264029 1961 264063 1989
rect 264091 1961 279237 1989
rect 279265 1961 279299 1989
rect 279327 1961 279361 1989
rect 279389 1961 279423 1989
rect 279451 1961 294597 1989
rect 294625 1961 294659 1989
rect 294687 1961 294721 1989
rect 294749 1961 294783 1989
rect 294811 1961 298248 1989
rect 298276 1961 298310 1989
rect 298338 1961 298372 1989
rect 298400 1961 298434 1989
rect 298462 1961 298990 1989
rect -958 1913 298990 1961
rect -478 -80 298510 -32
rect -478 -108 -430 -80
rect -402 -108 -368 -80
rect -340 -108 -306 -80
rect -278 -108 -244 -80
rect -216 -108 2757 -80
rect 2785 -108 2819 -80
rect 2847 -108 2881 -80
rect 2909 -108 2943 -80
rect 2971 -108 18117 -80
rect 18145 -108 18179 -80
rect 18207 -108 18241 -80
rect 18269 -108 18303 -80
rect 18331 -108 33477 -80
rect 33505 -108 33539 -80
rect 33567 -108 33601 -80
rect 33629 -108 33663 -80
rect 33691 -108 48837 -80
rect 48865 -108 48899 -80
rect 48927 -108 48961 -80
rect 48989 -108 49023 -80
rect 49051 -108 64197 -80
rect 64225 -108 64259 -80
rect 64287 -108 64321 -80
rect 64349 -108 64383 -80
rect 64411 -108 79557 -80
rect 79585 -108 79619 -80
rect 79647 -108 79681 -80
rect 79709 -108 79743 -80
rect 79771 -108 94917 -80
rect 94945 -108 94979 -80
rect 95007 -108 95041 -80
rect 95069 -108 95103 -80
rect 95131 -108 110277 -80
rect 110305 -108 110339 -80
rect 110367 -108 110401 -80
rect 110429 -108 110463 -80
rect 110491 -108 125637 -80
rect 125665 -108 125699 -80
rect 125727 -108 125761 -80
rect 125789 -108 125823 -80
rect 125851 -108 140997 -80
rect 141025 -108 141059 -80
rect 141087 -108 141121 -80
rect 141149 -108 141183 -80
rect 141211 -108 156357 -80
rect 156385 -108 156419 -80
rect 156447 -108 156481 -80
rect 156509 -108 156543 -80
rect 156571 -108 171717 -80
rect 171745 -108 171779 -80
rect 171807 -108 171841 -80
rect 171869 -108 171903 -80
rect 171931 -108 187077 -80
rect 187105 -108 187139 -80
rect 187167 -108 187201 -80
rect 187229 -108 187263 -80
rect 187291 -108 202437 -80
rect 202465 -108 202499 -80
rect 202527 -108 202561 -80
rect 202589 -108 202623 -80
rect 202651 -108 217797 -80
rect 217825 -108 217859 -80
rect 217887 -108 217921 -80
rect 217949 -108 217983 -80
rect 218011 -108 233157 -80
rect 233185 -108 233219 -80
rect 233247 -108 233281 -80
rect 233309 -108 233343 -80
rect 233371 -108 248517 -80
rect 248545 -108 248579 -80
rect 248607 -108 248641 -80
rect 248669 -108 248703 -80
rect 248731 -108 263877 -80
rect 263905 -108 263939 -80
rect 263967 -108 264001 -80
rect 264029 -108 264063 -80
rect 264091 -108 279237 -80
rect 279265 -108 279299 -80
rect 279327 -108 279361 -80
rect 279389 -108 279423 -80
rect 279451 -108 294597 -80
rect 294625 -108 294659 -80
rect 294687 -108 294721 -80
rect 294749 -108 294783 -80
rect 294811 -108 298248 -80
rect 298276 -108 298310 -80
rect 298338 -108 298372 -80
rect 298400 -108 298434 -80
rect 298462 -108 298510 -80
rect -478 -142 298510 -108
rect -478 -170 -430 -142
rect -402 -170 -368 -142
rect -340 -170 -306 -142
rect -278 -170 -244 -142
rect -216 -170 2757 -142
rect 2785 -170 2819 -142
rect 2847 -170 2881 -142
rect 2909 -170 2943 -142
rect 2971 -170 18117 -142
rect 18145 -170 18179 -142
rect 18207 -170 18241 -142
rect 18269 -170 18303 -142
rect 18331 -170 33477 -142
rect 33505 -170 33539 -142
rect 33567 -170 33601 -142
rect 33629 -170 33663 -142
rect 33691 -170 48837 -142
rect 48865 -170 48899 -142
rect 48927 -170 48961 -142
rect 48989 -170 49023 -142
rect 49051 -170 64197 -142
rect 64225 -170 64259 -142
rect 64287 -170 64321 -142
rect 64349 -170 64383 -142
rect 64411 -170 79557 -142
rect 79585 -170 79619 -142
rect 79647 -170 79681 -142
rect 79709 -170 79743 -142
rect 79771 -170 94917 -142
rect 94945 -170 94979 -142
rect 95007 -170 95041 -142
rect 95069 -170 95103 -142
rect 95131 -170 110277 -142
rect 110305 -170 110339 -142
rect 110367 -170 110401 -142
rect 110429 -170 110463 -142
rect 110491 -170 125637 -142
rect 125665 -170 125699 -142
rect 125727 -170 125761 -142
rect 125789 -170 125823 -142
rect 125851 -170 140997 -142
rect 141025 -170 141059 -142
rect 141087 -170 141121 -142
rect 141149 -170 141183 -142
rect 141211 -170 156357 -142
rect 156385 -170 156419 -142
rect 156447 -170 156481 -142
rect 156509 -170 156543 -142
rect 156571 -170 171717 -142
rect 171745 -170 171779 -142
rect 171807 -170 171841 -142
rect 171869 -170 171903 -142
rect 171931 -170 187077 -142
rect 187105 -170 187139 -142
rect 187167 -170 187201 -142
rect 187229 -170 187263 -142
rect 187291 -170 202437 -142
rect 202465 -170 202499 -142
rect 202527 -170 202561 -142
rect 202589 -170 202623 -142
rect 202651 -170 217797 -142
rect 217825 -170 217859 -142
rect 217887 -170 217921 -142
rect 217949 -170 217983 -142
rect 218011 -170 233157 -142
rect 233185 -170 233219 -142
rect 233247 -170 233281 -142
rect 233309 -170 233343 -142
rect 233371 -170 248517 -142
rect 248545 -170 248579 -142
rect 248607 -170 248641 -142
rect 248669 -170 248703 -142
rect 248731 -170 263877 -142
rect 263905 -170 263939 -142
rect 263967 -170 264001 -142
rect 264029 -170 264063 -142
rect 264091 -170 279237 -142
rect 279265 -170 279299 -142
rect 279327 -170 279361 -142
rect 279389 -170 279423 -142
rect 279451 -170 294597 -142
rect 294625 -170 294659 -142
rect 294687 -170 294721 -142
rect 294749 -170 294783 -142
rect 294811 -170 298248 -142
rect 298276 -170 298310 -142
rect 298338 -170 298372 -142
rect 298400 -170 298434 -142
rect 298462 -170 298510 -142
rect -478 -204 298510 -170
rect -478 -232 -430 -204
rect -402 -232 -368 -204
rect -340 -232 -306 -204
rect -278 -232 -244 -204
rect -216 -232 2757 -204
rect 2785 -232 2819 -204
rect 2847 -232 2881 -204
rect 2909 -232 2943 -204
rect 2971 -232 18117 -204
rect 18145 -232 18179 -204
rect 18207 -232 18241 -204
rect 18269 -232 18303 -204
rect 18331 -232 33477 -204
rect 33505 -232 33539 -204
rect 33567 -232 33601 -204
rect 33629 -232 33663 -204
rect 33691 -232 48837 -204
rect 48865 -232 48899 -204
rect 48927 -232 48961 -204
rect 48989 -232 49023 -204
rect 49051 -232 64197 -204
rect 64225 -232 64259 -204
rect 64287 -232 64321 -204
rect 64349 -232 64383 -204
rect 64411 -232 79557 -204
rect 79585 -232 79619 -204
rect 79647 -232 79681 -204
rect 79709 -232 79743 -204
rect 79771 -232 94917 -204
rect 94945 -232 94979 -204
rect 95007 -232 95041 -204
rect 95069 -232 95103 -204
rect 95131 -232 110277 -204
rect 110305 -232 110339 -204
rect 110367 -232 110401 -204
rect 110429 -232 110463 -204
rect 110491 -232 125637 -204
rect 125665 -232 125699 -204
rect 125727 -232 125761 -204
rect 125789 -232 125823 -204
rect 125851 -232 140997 -204
rect 141025 -232 141059 -204
rect 141087 -232 141121 -204
rect 141149 -232 141183 -204
rect 141211 -232 156357 -204
rect 156385 -232 156419 -204
rect 156447 -232 156481 -204
rect 156509 -232 156543 -204
rect 156571 -232 171717 -204
rect 171745 -232 171779 -204
rect 171807 -232 171841 -204
rect 171869 -232 171903 -204
rect 171931 -232 187077 -204
rect 187105 -232 187139 -204
rect 187167 -232 187201 -204
rect 187229 -232 187263 -204
rect 187291 -232 202437 -204
rect 202465 -232 202499 -204
rect 202527 -232 202561 -204
rect 202589 -232 202623 -204
rect 202651 -232 217797 -204
rect 217825 -232 217859 -204
rect 217887 -232 217921 -204
rect 217949 -232 217983 -204
rect 218011 -232 233157 -204
rect 233185 -232 233219 -204
rect 233247 -232 233281 -204
rect 233309 -232 233343 -204
rect 233371 -232 248517 -204
rect 248545 -232 248579 -204
rect 248607 -232 248641 -204
rect 248669 -232 248703 -204
rect 248731 -232 263877 -204
rect 263905 -232 263939 -204
rect 263967 -232 264001 -204
rect 264029 -232 264063 -204
rect 264091 -232 279237 -204
rect 279265 -232 279299 -204
rect 279327 -232 279361 -204
rect 279389 -232 279423 -204
rect 279451 -232 294597 -204
rect 294625 -232 294659 -204
rect 294687 -232 294721 -204
rect 294749 -232 294783 -204
rect 294811 -232 298248 -204
rect 298276 -232 298310 -204
rect 298338 -232 298372 -204
rect 298400 -232 298434 -204
rect 298462 -232 298510 -204
rect -478 -266 298510 -232
rect -478 -294 -430 -266
rect -402 -294 -368 -266
rect -340 -294 -306 -266
rect -278 -294 -244 -266
rect -216 -294 2757 -266
rect 2785 -294 2819 -266
rect 2847 -294 2881 -266
rect 2909 -294 2943 -266
rect 2971 -294 18117 -266
rect 18145 -294 18179 -266
rect 18207 -294 18241 -266
rect 18269 -294 18303 -266
rect 18331 -294 33477 -266
rect 33505 -294 33539 -266
rect 33567 -294 33601 -266
rect 33629 -294 33663 -266
rect 33691 -294 48837 -266
rect 48865 -294 48899 -266
rect 48927 -294 48961 -266
rect 48989 -294 49023 -266
rect 49051 -294 64197 -266
rect 64225 -294 64259 -266
rect 64287 -294 64321 -266
rect 64349 -294 64383 -266
rect 64411 -294 79557 -266
rect 79585 -294 79619 -266
rect 79647 -294 79681 -266
rect 79709 -294 79743 -266
rect 79771 -294 94917 -266
rect 94945 -294 94979 -266
rect 95007 -294 95041 -266
rect 95069 -294 95103 -266
rect 95131 -294 110277 -266
rect 110305 -294 110339 -266
rect 110367 -294 110401 -266
rect 110429 -294 110463 -266
rect 110491 -294 125637 -266
rect 125665 -294 125699 -266
rect 125727 -294 125761 -266
rect 125789 -294 125823 -266
rect 125851 -294 140997 -266
rect 141025 -294 141059 -266
rect 141087 -294 141121 -266
rect 141149 -294 141183 -266
rect 141211 -294 156357 -266
rect 156385 -294 156419 -266
rect 156447 -294 156481 -266
rect 156509 -294 156543 -266
rect 156571 -294 171717 -266
rect 171745 -294 171779 -266
rect 171807 -294 171841 -266
rect 171869 -294 171903 -266
rect 171931 -294 187077 -266
rect 187105 -294 187139 -266
rect 187167 -294 187201 -266
rect 187229 -294 187263 -266
rect 187291 -294 202437 -266
rect 202465 -294 202499 -266
rect 202527 -294 202561 -266
rect 202589 -294 202623 -266
rect 202651 -294 217797 -266
rect 217825 -294 217859 -266
rect 217887 -294 217921 -266
rect 217949 -294 217983 -266
rect 218011 -294 233157 -266
rect 233185 -294 233219 -266
rect 233247 -294 233281 -266
rect 233309 -294 233343 -266
rect 233371 -294 248517 -266
rect 248545 -294 248579 -266
rect 248607 -294 248641 -266
rect 248669 -294 248703 -266
rect 248731 -294 263877 -266
rect 263905 -294 263939 -266
rect 263967 -294 264001 -266
rect 264029 -294 264063 -266
rect 264091 -294 279237 -266
rect 279265 -294 279299 -266
rect 279327 -294 279361 -266
rect 279389 -294 279423 -266
rect 279451 -294 294597 -266
rect 294625 -294 294659 -266
rect 294687 -294 294721 -266
rect 294749 -294 294783 -266
rect 294811 -294 298248 -266
rect 298276 -294 298310 -266
rect 298338 -294 298372 -266
rect 298400 -294 298434 -266
rect 298462 -294 298510 -266
rect -478 -342 298510 -294
rect -958 -560 298990 -512
rect -958 -588 -910 -560
rect -882 -588 -848 -560
rect -820 -588 -786 -560
rect -758 -588 -724 -560
rect -696 -588 4617 -560
rect 4645 -588 4679 -560
rect 4707 -588 4741 -560
rect 4769 -588 4803 -560
rect 4831 -588 19977 -560
rect 20005 -588 20039 -560
rect 20067 -588 20101 -560
rect 20129 -588 20163 -560
rect 20191 -588 35337 -560
rect 35365 -588 35399 -560
rect 35427 -588 35461 -560
rect 35489 -588 35523 -560
rect 35551 -588 50697 -560
rect 50725 -588 50759 -560
rect 50787 -588 50821 -560
rect 50849 -588 50883 -560
rect 50911 -588 66057 -560
rect 66085 -588 66119 -560
rect 66147 -588 66181 -560
rect 66209 -588 66243 -560
rect 66271 -588 81417 -560
rect 81445 -588 81479 -560
rect 81507 -588 81541 -560
rect 81569 -588 81603 -560
rect 81631 -588 96777 -560
rect 96805 -588 96839 -560
rect 96867 -588 96901 -560
rect 96929 -588 96963 -560
rect 96991 -588 112137 -560
rect 112165 -588 112199 -560
rect 112227 -588 112261 -560
rect 112289 -588 112323 -560
rect 112351 -588 127497 -560
rect 127525 -588 127559 -560
rect 127587 -588 127621 -560
rect 127649 -588 127683 -560
rect 127711 -588 142857 -560
rect 142885 -588 142919 -560
rect 142947 -588 142981 -560
rect 143009 -588 143043 -560
rect 143071 -588 158217 -560
rect 158245 -588 158279 -560
rect 158307 -588 158341 -560
rect 158369 -588 158403 -560
rect 158431 -588 173577 -560
rect 173605 -588 173639 -560
rect 173667 -588 173701 -560
rect 173729 -588 173763 -560
rect 173791 -588 188937 -560
rect 188965 -588 188999 -560
rect 189027 -588 189061 -560
rect 189089 -588 189123 -560
rect 189151 -588 204297 -560
rect 204325 -588 204359 -560
rect 204387 -588 204421 -560
rect 204449 -588 204483 -560
rect 204511 -588 219657 -560
rect 219685 -588 219719 -560
rect 219747 -588 219781 -560
rect 219809 -588 219843 -560
rect 219871 -588 235017 -560
rect 235045 -588 235079 -560
rect 235107 -588 235141 -560
rect 235169 -588 235203 -560
rect 235231 -588 250377 -560
rect 250405 -588 250439 -560
rect 250467 -588 250501 -560
rect 250529 -588 250563 -560
rect 250591 -588 265737 -560
rect 265765 -588 265799 -560
rect 265827 -588 265861 -560
rect 265889 -588 265923 -560
rect 265951 -588 281097 -560
rect 281125 -588 281159 -560
rect 281187 -588 281221 -560
rect 281249 -588 281283 -560
rect 281311 -588 296457 -560
rect 296485 -588 296519 -560
rect 296547 -588 296581 -560
rect 296609 -588 296643 -560
rect 296671 -588 298728 -560
rect 298756 -588 298790 -560
rect 298818 -588 298852 -560
rect 298880 -588 298914 -560
rect 298942 -588 298990 -560
rect -958 -622 298990 -588
rect -958 -650 -910 -622
rect -882 -650 -848 -622
rect -820 -650 -786 -622
rect -758 -650 -724 -622
rect -696 -650 4617 -622
rect 4645 -650 4679 -622
rect 4707 -650 4741 -622
rect 4769 -650 4803 -622
rect 4831 -650 19977 -622
rect 20005 -650 20039 -622
rect 20067 -650 20101 -622
rect 20129 -650 20163 -622
rect 20191 -650 35337 -622
rect 35365 -650 35399 -622
rect 35427 -650 35461 -622
rect 35489 -650 35523 -622
rect 35551 -650 50697 -622
rect 50725 -650 50759 -622
rect 50787 -650 50821 -622
rect 50849 -650 50883 -622
rect 50911 -650 66057 -622
rect 66085 -650 66119 -622
rect 66147 -650 66181 -622
rect 66209 -650 66243 -622
rect 66271 -650 81417 -622
rect 81445 -650 81479 -622
rect 81507 -650 81541 -622
rect 81569 -650 81603 -622
rect 81631 -650 96777 -622
rect 96805 -650 96839 -622
rect 96867 -650 96901 -622
rect 96929 -650 96963 -622
rect 96991 -650 112137 -622
rect 112165 -650 112199 -622
rect 112227 -650 112261 -622
rect 112289 -650 112323 -622
rect 112351 -650 127497 -622
rect 127525 -650 127559 -622
rect 127587 -650 127621 -622
rect 127649 -650 127683 -622
rect 127711 -650 142857 -622
rect 142885 -650 142919 -622
rect 142947 -650 142981 -622
rect 143009 -650 143043 -622
rect 143071 -650 158217 -622
rect 158245 -650 158279 -622
rect 158307 -650 158341 -622
rect 158369 -650 158403 -622
rect 158431 -650 173577 -622
rect 173605 -650 173639 -622
rect 173667 -650 173701 -622
rect 173729 -650 173763 -622
rect 173791 -650 188937 -622
rect 188965 -650 188999 -622
rect 189027 -650 189061 -622
rect 189089 -650 189123 -622
rect 189151 -650 204297 -622
rect 204325 -650 204359 -622
rect 204387 -650 204421 -622
rect 204449 -650 204483 -622
rect 204511 -650 219657 -622
rect 219685 -650 219719 -622
rect 219747 -650 219781 -622
rect 219809 -650 219843 -622
rect 219871 -650 235017 -622
rect 235045 -650 235079 -622
rect 235107 -650 235141 -622
rect 235169 -650 235203 -622
rect 235231 -650 250377 -622
rect 250405 -650 250439 -622
rect 250467 -650 250501 -622
rect 250529 -650 250563 -622
rect 250591 -650 265737 -622
rect 265765 -650 265799 -622
rect 265827 -650 265861 -622
rect 265889 -650 265923 -622
rect 265951 -650 281097 -622
rect 281125 -650 281159 -622
rect 281187 -650 281221 -622
rect 281249 -650 281283 -622
rect 281311 -650 296457 -622
rect 296485 -650 296519 -622
rect 296547 -650 296581 -622
rect 296609 -650 296643 -622
rect 296671 -650 298728 -622
rect 298756 -650 298790 -622
rect 298818 -650 298852 -622
rect 298880 -650 298914 -622
rect 298942 -650 298990 -622
rect -958 -684 298990 -650
rect -958 -712 -910 -684
rect -882 -712 -848 -684
rect -820 -712 -786 -684
rect -758 -712 -724 -684
rect -696 -712 4617 -684
rect 4645 -712 4679 -684
rect 4707 -712 4741 -684
rect 4769 -712 4803 -684
rect 4831 -712 19977 -684
rect 20005 -712 20039 -684
rect 20067 -712 20101 -684
rect 20129 -712 20163 -684
rect 20191 -712 35337 -684
rect 35365 -712 35399 -684
rect 35427 -712 35461 -684
rect 35489 -712 35523 -684
rect 35551 -712 50697 -684
rect 50725 -712 50759 -684
rect 50787 -712 50821 -684
rect 50849 -712 50883 -684
rect 50911 -712 66057 -684
rect 66085 -712 66119 -684
rect 66147 -712 66181 -684
rect 66209 -712 66243 -684
rect 66271 -712 81417 -684
rect 81445 -712 81479 -684
rect 81507 -712 81541 -684
rect 81569 -712 81603 -684
rect 81631 -712 96777 -684
rect 96805 -712 96839 -684
rect 96867 -712 96901 -684
rect 96929 -712 96963 -684
rect 96991 -712 112137 -684
rect 112165 -712 112199 -684
rect 112227 -712 112261 -684
rect 112289 -712 112323 -684
rect 112351 -712 127497 -684
rect 127525 -712 127559 -684
rect 127587 -712 127621 -684
rect 127649 -712 127683 -684
rect 127711 -712 142857 -684
rect 142885 -712 142919 -684
rect 142947 -712 142981 -684
rect 143009 -712 143043 -684
rect 143071 -712 158217 -684
rect 158245 -712 158279 -684
rect 158307 -712 158341 -684
rect 158369 -712 158403 -684
rect 158431 -712 173577 -684
rect 173605 -712 173639 -684
rect 173667 -712 173701 -684
rect 173729 -712 173763 -684
rect 173791 -712 188937 -684
rect 188965 -712 188999 -684
rect 189027 -712 189061 -684
rect 189089 -712 189123 -684
rect 189151 -712 204297 -684
rect 204325 -712 204359 -684
rect 204387 -712 204421 -684
rect 204449 -712 204483 -684
rect 204511 -712 219657 -684
rect 219685 -712 219719 -684
rect 219747 -712 219781 -684
rect 219809 -712 219843 -684
rect 219871 -712 235017 -684
rect 235045 -712 235079 -684
rect 235107 -712 235141 -684
rect 235169 -712 235203 -684
rect 235231 -712 250377 -684
rect 250405 -712 250439 -684
rect 250467 -712 250501 -684
rect 250529 -712 250563 -684
rect 250591 -712 265737 -684
rect 265765 -712 265799 -684
rect 265827 -712 265861 -684
rect 265889 -712 265923 -684
rect 265951 -712 281097 -684
rect 281125 -712 281159 -684
rect 281187 -712 281221 -684
rect 281249 -712 281283 -684
rect 281311 -712 296457 -684
rect 296485 -712 296519 -684
rect 296547 -712 296581 -684
rect 296609 -712 296643 -684
rect 296671 -712 298728 -684
rect 298756 -712 298790 -684
rect 298818 -712 298852 -684
rect 298880 -712 298914 -684
rect 298942 -712 298990 -684
rect -958 -746 298990 -712
rect -958 -774 -910 -746
rect -882 -774 -848 -746
rect -820 -774 -786 -746
rect -758 -774 -724 -746
rect -696 -774 4617 -746
rect 4645 -774 4679 -746
rect 4707 -774 4741 -746
rect 4769 -774 4803 -746
rect 4831 -774 19977 -746
rect 20005 -774 20039 -746
rect 20067 -774 20101 -746
rect 20129 -774 20163 -746
rect 20191 -774 35337 -746
rect 35365 -774 35399 -746
rect 35427 -774 35461 -746
rect 35489 -774 35523 -746
rect 35551 -774 50697 -746
rect 50725 -774 50759 -746
rect 50787 -774 50821 -746
rect 50849 -774 50883 -746
rect 50911 -774 66057 -746
rect 66085 -774 66119 -746
rect 66147 -774 66181 -746
rect 66209 -774 66243 -746
rect 66271 -774 81417 -746
rect 81445 -774 81479 -746
rect 81507 -774 81541 -746
rect 81569 -774 81603 -746
rect 81631 -774 96777 -746
rect 96805 -774 96839 -746
rect 96867 -774 96901 -746
rect 96929 -774 96963 -746
rect 96991 -774 112137 -746
rect 112165 -774 112199 -746
rect 112227 -774 112261 -746
rect 112289 -774 112323 -746
rect 112351 -774 127497 -746
rect 127525 -774 127559 -746
rect 127587 -774 127621 -746
rect 127649 -774 127683 -746
rect 127711 -774 142857 -746
rect 142885 -774 142919 -746
rect 142947 -774 142981 -746
rect 143009 -774 143043 -746
rect 143071 -774 158217 -746
rect 158245 -774 158279 -746
rect 158307 -774 158341 -746
rect 158369 -774 158403 -746
rect 158431 -774 173577 -746
rect 173605 -774 173639 -746
rect 173667 -774 173701 -746
rect 173729 -774 173763 -746
rect 173791 -774 188937 -746
rect 188965 -774 188999 -746
rect 189027 -774 189061 -746
rect 189089 -774 189123 -746
rect 189151 -774 204297 -746
rect 204325 -774 204359 -746
rect 204387 -774 204421 -746
rect 204449 -774 204483 -746
rect 204511 -774 219657 -746
rect 219685 -774 219719 -746
rect 219747 -774 219781 -746
rect 219809 -774 219843 -746
rect 219871 -774 235017 -746
rect 235045 -774 235079 -746
rect 235107 -774 235141 -746
rect 235169 -774 235203 -746
rect 235231 -774 250377 -746
rect 250405 -774 250439 -746
rect 250467 -774 250501 -746
rect 250529 -774 250563 -746
rect 250591 -774 265737 -746
rect 265765 -774 265799 -746
rect 265827 -774 265861 -746
rect 265889 -774 265923 -746
rect 265951 -774 281097 -746
rect 281125 -774 281159 -746
rect 281187 -774 281221 -746
rect 281249 -774 281283 -746
rect 281311 -774 296457 -746
rect 296485 -774 296519 -746
rect 296547 -774 296581 -746
rect 296609 -774 296643 -746
rect 296671 -774 298728 -746
rect 298756 -774 298790 -746
rect 298818 -774 298852 -746
rect 298880 -774 298914 -746
rect 298942 -774 298990 -746
rect -958 -822 298990 -774
use top_design_mux  top_design_mux
timestamp 0
transform 1 0 30000 0 1 130000
box 0 0 240000 30000
use top_raybox_zero_fsm  top_raybox_zero_fsm
timestamp 0
transform 1 0 20000 0 1 170000
box 513 0 65856 99206
use top_raybox_zero_fsm  top_raybox_zero_fsm2
timestamp 0
transform 1 0 100000 0 1 170000
box 513 0 65856 99206
use top_solo_squash  top_solo_squash
timestamp 0
transform 1 0 235000 0 1 170000
box 629 0 20035 20819
use top_vga_spi_rom  top_vga_spi_rom
timestamp 0
transform 1 0 180000 0 1 170000
box 629 0 24403 25191
use urish_simon_says  urish_simon_says
timestamp 0
transform 1 0 100000 0 1 95000
box 629 1525 29331 30000
use user_proj_cpu  user_proj_cpu
timestamp 0
transform 1 0 160000 0 1 7000
box 629 401 115571 118024
use wrapped_wb_hyperram  wrapped_wb_hyperram
timestamp 0
transform 1 0 14000 0 1 75000
box 629 0 79339 30000
<< labels >>
flabel metal3 s 297780 3556 298500 3668 0 FreeSans 448 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 297780 201796 298500 201908 0 FreeSans 448 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 297780 221620 298500 221732 0 FreeSans 448 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 297780 241444 298500 241556 0 FreeSans 448 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 297780 261268 298500 261380 0 FreeSans 448 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 297780 281092 298500 281204 0 FreeSans 448 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 292348 297780 292460 298500 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 259252 297780 259364 298500 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 226156 297780 226268 298500 0 FreeSans 448 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 193060 297780 193172 298500 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 159964 297780 160076 298500 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 297780 23380 298500 23492 0 FreeSans 448 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 126868 297780 126980 298500 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 93772 297780 93884 298500 0 FreeSans 448 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 60676 297780 60788 298500 0 FreeSans 448 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 27580 297780 27692 298500 0 FreeSans 448 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -480 293580 240 293692 0 FreeSans 448 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -480 272412 240 272524 0 FreeSans 448 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -480 251244 240 251356 0 FreeSans 448 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -480 230076 240 230188 0 FreeSans 448 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -480 208908 240 209020 0 FreeSans 448 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -480 187740 240 187852 0 FreeSans 448 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 297780 43204 298500 43316 0 FreeSans 448 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -480 166572 240 166684 0 FreeSans 448 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -480 145404 240 145516 0 FreeSans 448 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -480 124236 240 124348 0 FreeSans 448 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -480 103068 240 103180 0 FreeSans 448 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -480 81900 240 82012 0 FreeSans 448 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -480 60732 240 60844 0 FreeSans 448 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -480 39564 240 39676 0 FreeSans 448 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -480 18396 240 18508 0 FreeSans 448 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 297780 63028 298500 63140 0 FreeSans 448 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 297780 82852 298500 82964 0 FreeSans 448 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 297780 102676 298500 102788 0 FreeSans 448 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 297780 122500 298500 122612 0 FreeSans 448 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 297780 142324 298500 142436 0 FreeSans 448 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 297780 162148 298500 162260 0 FreeSans 448 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 297780 181972 298500 182084 0 FreeSans 448 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 297780 16772 298500 16884 0 FreeSans 448 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 297780 215012 298500 215124 0 FreeSans 448 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 297780 234836 298500 234948 0 FreeSans 448 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 297780 254660 298500 254772 0 FreeSans 448 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 297780 274484 298500 274596 0 FreeSans 448 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 297780 294308 298500 294420 0 FreeSans 448 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 270284 297780 270396 298500 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 237188 297780 237300 298500 0 FreeSans 448 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 204092 297780 204204 298500 0 FreeSans 448 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 170996 297780 171108 298500 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 137900 297780 138012 298500 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 297780 36596 298500 36708 0 FreeSans 448 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 104804 297780 104916 298500 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 71708 297780 71820 298500 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 38612 297780 38724 298500 0 FreeSans 448 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 5516 297780 5628 298500 0 FreeSans 448 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -480 279468 240 279580 0 FreeSans 448 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -480 258300 240 258412 0 FreeSans 448 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -480 237132 240 237244 0 FreeSans 448 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -480 215964 240 216076 0 FreeSans 448 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -480 194796 240 194908 0 FreeSans 448 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -480 173628 240 173740 0 FreeSans 448 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 297780 56420 298500 56532 0 FreeSans 448 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -480 152460 240 152572 0 FreeSans 448 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -480 131292 240 131404 0 FreeSans 448 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -480 110124 240 110236 0 FreeSans 448 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -480 88956 240 89068 0 FreeSans 448 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -480 67788 240 67900 0 FreeSans 448 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -480 46620 240 46732 0 FreeSans 448 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -480 25452 240 25564 0 FreeSans 448 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -480 4284 240 4396 0 FreeSans 448 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 297780 76244 298500 76356 0 FreeSans 448 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 297780 96068 298500 96180 0 FreeSans 448 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 297780 115892 298500 116004 0 FreeSans 448 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 297780 135716 298500 135828 0 FreeSans 448 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 297780 155540 298500 155652 0 FreeSans 448 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 297780 175364 298500 175476 0 FreeSans 448 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 297780 195188 298500 195300 0 FreeSans 448 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 297780 10164 298500 10276 0 FreeSans 448 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 297780 208404 298500 208516 0 FreeSans 448 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 297780 228228 298500 228340 0 FreeSans 448 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 297780 248052 298500 248164 0 FreeSans 448 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 297780 267876 298500 267988 0 FreeSans 448 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 297780 287700 298500 287812 0 FreeSans 448 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 281316 297780 281428 298500 0 FreeSans 448 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 248220 297780 248332 298500 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 215124 297780 215236 298500 0 FreeSans 448 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 182028 297780 182140 298500 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 148932 297780 149044 298500 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 297780 29988 298500 30100 0 FreeSans 448 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 115836 297780 115948 298500 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 82740 297780 82852 298500 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 49644 297780 49756 298500 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 16548 297780 16660 298500 0 FreeSans 448 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -480 286524 240 286636 0 FreeSans 448 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -480 265356 240 265468 0 FreeSans 448 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -480 244188 240 244300 0 FreeSans 448 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -480 223020 240 223132 0 FreeSans 448 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -480 201852 240 201964 0 FreeSans 448 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -480 180684 240 180796 0 FreeSans 448 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 297780 49812 298500 49924 0 FreeSans 448 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -480 159516 240 159628 0 FreeSans 448 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -480 138348 240 138460 0 FreeSans 448 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -480 117180 240 117292 0 FreeSans 448 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -480 96012 240 96124 0 FreeSans 448 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -480 74844 240 74956 0 FreeSans 448 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -480 53676 240 53788 0 FreeSans 448 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -480 32508 240 32620 0 FreeSans 448 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -480 11340 240 11452 0 FreeSans 448 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 297780 69636 298500 69748 0 FreeSans 448 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 297780 89460 298500 89572 0 FreeSans 448 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 297780 109284 298500 109396 0 FreeSans 448 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 297780 129108 298500 129220 0 FreeSans 448 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 297780 148932 298500 149044 0 FreeSans 448 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 297780 168756 298500 168868 0 FreeSans 448 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 297780 188580 298500 188692 0 FreeSans 448 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 106596 -480 106708 240 0 FreeSans 448 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 135156 -480 135268 240 0 FreeSans 448 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 138012 -480 138124 240 0 FreeSans 448 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 140868 -480 140980 240 0 FreeSans 448 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 143724 -480 143836 240 0 FreeSans 448 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 146580 -480 146692 240 0 FreeSans 448 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 149436 -480 149548 240 0 FreeSans 448 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 152292 -480 152404 240 0 FreeSans 448 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 155148 -480 155260 240 0 FreeSans 448 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 158004 -480 158116 240 0 FreeSans 448 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 160860 -480 160972 240 0 FreeSans 448 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 109452 -480 109564 240 0 FreeSans 448 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 163716 -480 163828 240 0 FreeSans 448 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 166572 -480 166684 240 0 FreeSans 448 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 169428 -480 169540 240 0 FreeSans 448 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 172284 -480 172396 240 0 FreeSans 448 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 175140 -480 175252 240 0 FreeSans 448 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 177996 -480 178108 240 0 FreeSans 448 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 180852 -480 180964 240 0 FreeSans 448 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 183708 -480 183820 240 0 FreeSans 448 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 186564 -480 186676 240 0 FreeSans 448 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 189420 -480 189532 240 0 FreeSans 448 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 112308 -480 112420 240 0 FreeSans 448 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 192276 -480 192388 240 0 FreeSans 448 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 195132 -480 195244 240 0 FreeSans 448 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 197988 -480 198100 240 0 FreeSans 448 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 200844 -480 200956 240 0 FreeSans 448 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 203700 -480 203812 240 0 FreeSans 448 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 206556 -480 206668 240 0 FreeSans 448 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 209412 -480 209524 240 0 FreeSans 448 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 212268 -480 212380 240 0 FreeSans 448 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 215124 -480 215236 240 0 FreeSans 448 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 217980 -480 218092 240 0 FreeSans 448 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 115164 -480 115276 240 0 FreeSans 448 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 220836 -480 220948 240 0 FreeSans 448 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 223692 -480 223804 240 0 FreeSans 448 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 226548 -480 226660 240 0 FreeSans 448 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 229404 -480 229516 240 0 FreeSans 448 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 232260 -480 232372 240 0 FreeSans 448 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 235116 -480 235228 240 0 FreeSans 448 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 237972 -480 238084 240 0 FreeSans 448 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 240828 -480 240940 240 0 FreeSans 448 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 243684 -480 243796 240 0 FreeSans 448 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 246540 -480 246652 240 0 FreeSans 448 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 118020 -480 118132 240 0 FreeSans 448 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 249396 -480 249508 240 0 FreeSans 448 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 252252 -480 252364 240 0 FreeSans 448 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 255108 -480 255220 240 0 FreeSans 448 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 257964 -480 258076 240 0 FreeSans 448 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 260820 -480 260932 240 0 FreeSans 448 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 263676 -480 263788 240 0 FreeSans 448 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 266532 -480 266644 240 0 FreeSans 448 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 269388 -480 269500 240 0 FreeSans 448 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 272244 -480 272356 240 0 FreeSans 448 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 275100 -480 275212 240 0 FreeSans 448 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 120876 -480 120988 240 0 FreeSans 448 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 277956 -480 278068 240 0 FreeSans 448 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 280812 -480 280924 240 0 FreeSans 448 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 283668 -480 283780 240 0 FreeSans 448 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 286524 -480 286636 240 0 FreeSans 448 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 123732 -480 123844 240 0 FreeSans 448 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 126588 -480 126700 240 0 FreeSans 448 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 129444 -480 129556 240 0 FreeSans 448 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 132300 -480 132412 240 0 FreeSans 448 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 107548 -480 107660 240 0 FreeSans 448 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 136108 -480 136220 240 0 FreeSans 448 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 138964 -480 139076 240 0 FreeSans 448 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 141820 -480 141932 240 0 FreeSans 448 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 144676 -480 144788 240 0 FreeSans 448 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 147532 -480 147644 240 0 FreeSans 448 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 150388 -480 150500 240 0 FreeSans 448 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 153244 -480 153356 240 0 FreeSans 448 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 156100 -480 156212 240 0 FreeSans 448 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 158956 -480 159068 240 0 FreeSans 448 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 161812 -480 161924 240 0 FreeSans 448 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 110404 -480 110516 240 0 FreeSans 448 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 164668 -480 164780 240 0 FreeSans 448 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 167524 -480 167636 240 0 FreeSans 448 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 170380 -480 170492 240 0 FreeSans 448 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 173236 -480 173348 240 0 FreeSans 448 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 176092 -480 176204 240 0 FreeSans 448 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 178948 -480 179060 240 0 FreeSans 448 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 181804 -480 181916 240 0 FreeSans 448 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 184660 -480 184772 240 0 FreeSans 448 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 187516 -480 187628 240 0 FreeSans 448 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 190372 -480 190484 240 0 FreeSans 448 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 113260 -480 113372 240 0 FreeSans 448 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 193228 -480 193340 240 0 FreeSans 448 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 196084 -480 196196 240 0 FreeSans 448 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 198940 -480 199052 240 0 FreeSans 448 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 201796 -480 201908 240 0 FreeSans 448 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 204652 -480 204764 240 0 FreeSans 448 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 207508 -480 207620 240 0 FreeSans 448 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 210364 -480 210476 240 0 FreeSans 448 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 213220 -480 213332 240 0 FreeSans 448 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 216076 -480 216188 240 0 FreeSans 448 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 218932 -480 219044 240 0 FreeSans 448 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 116116 -480 116228 240 0 FreeSans 448 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 221788 -480 221900 240 0 FreeSans 448 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 224644 -480 224756 240 0 FreeSans 448 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 227500 -480 227612 240 0 FreeSans 448 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 230356 -480 230468 240 0 FreeSans 448 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 233212 -480 233324 240 0 FreeSans 448 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 236068 -480 236180 240 0 FreeSans 448 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 238924 -480 239036 240 0 FreeSans 448 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 241780 -480 241892 240 0 FreeSans 448 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 244636 -480 244748 240 0 FreeSans 448 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 247492 -480 247604 240 0 FreeSans 448 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 118972 -480 119084 240 0 FreeSans 448 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 250348 -480 250460 240 0 FreeSans 448 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 253204 -480 253316 240 0 FreeSans 448 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 256060 -480 256172 240 0 FreeSans 448 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 258916 -480 259028 240 0 FreeSans 448 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 261772 -480 261884 240 0 FreeSans 448 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 264628 -480 264740 240 0 FreeSans 448 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 267484 -480 267596 240 0 FreeSans 448 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 270340 -480 270452 240 0 FreeSans 448 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 273196 -480 273308 240 0 FreeSans 448 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 276052 -480 276164 240 0 FreeSans 448 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 121828 -480 121940 240 0 FreeSans 448 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 278908 -480 279020 240 0 FreeSans 448 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 281764 -480 281876 240 0 FreeSans 448 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 284620 -480 284732 240 0 FreeSans 448 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 287476 -480 287588 240 0 FreeSans 448 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 124684 -480 124796 240 0 FreeSans 448 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 127540 -480 127652 240 0 FreeSans 448 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 130396 -480 130508 240 0 FreeSans 448 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 133252 -480 133364 240 0 FreeSans 448 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 108500 -480 108612 240 0 FreeSans 448 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 137060 -480 137172 240 0 FreeSans 448 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 139916 -480 140028 240 0 FreeSans 448 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 142772 -480 142884 240 0 FreeSans 448 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 145628 -480 145740 240 0 FreeSans 448 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 148484 -480 148596 240 0 FreeSans 448 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 151340 -480 151452 240 0 FreeSans 448 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 154196 -480 154308 240 0 FreeSans 448 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 157052 -480 157164 240 0 FreeSans 448 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 159908 -480 160020 240 0 FreeSans 448 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 162764 -480 162876 240 0 FreeSans 448 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 111356 -480 111468 240 0 FreeSans 448 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 165620 -480 165732 240 0 FreeSans 448 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 168476 -480 168588 240 0 FreeSans 448 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 171332 -480 171444 240 0 FreeSans 448 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 174188 -480 174300 240 0 FreeSans 448 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 177044 -480 177156 240 0 FreeSans 448 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 179900 -480 180012 240 0 FreeSans 448 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 182756 -480 182868 240 0 FreeSans 448 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 185612 -480 185724 240 0 FreeSans 448 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 188468 -480 188580 240 0 FreeSans 448 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 191324 -480 191436 240 0 FreeSans 448 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 114212 -480 114324 240 0 FreeSans 448 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 194180 -480 194292 240 0 FreeSans 448 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 197036 -480 197148 240 0 FreeSans 448 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 199892 -480 200004 240 0 FreeSans 448 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 202748 -480 202860 240 0 FreeSans 448 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 205604 -480 205716 240 0 FreeSans 448 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 208460 -480 208572 240 0 FreeSans 448 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 211316 -480 211428 240 0 FreeSans 448 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 214172 -480 214284 240 0 FreeSans 448 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 217028 -480 217140 240 0 FreeSans 448 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 219884 -480 219996 240 0 FreeSans 448 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 117068 -480 117180 240 0 FreeSans 448 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 222740 -480 222852 240 0 FreeSans 448 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 225596 -480 225708 240 0 FreeSans 448 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 228452 -480 228564 240 0 FreeSans 448 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 231308 -480 231420 240 0 FreeSans 448 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 234164 -480 234276 240 0 FreeSans 448 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 237020 -480 237132 240 0 FreeSans 448 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 239876 -480 239988 240 0 FreeSans 448 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 242732 -480 242844 240 0 FreeSans 448 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 245588 -480 245700 240 0 FreeSans 448 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 248444 -480 248556 240 0 FreeSans 448 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 119924 -480 120036 240 0 FreeSans 448 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 251300 -480 251412 240 0 FreeSans 448 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 254156 -480 254268 240 0 FreeSans 448 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 257012 -480 257124 240 0 FreeSans 448 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 259868 -480 259980 240 0 FreeSans 448 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 262724 -480 262836 240 0 FreeSans 448 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 265580 -480 265692 240 0 FreeSans 448 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 268436 -480 268548 240 0 FreeSans 448 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 271292 -480 271404 240 0 FreeSans 448 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 274148 -480 274260 240 0 FreeSans 448 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 277004 -480 277116 240 0 FreeSans 448 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 122780 -480 122892 240 0 FreeSans 448 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 279860 -480 279972 240 0 FreeSans 448 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 282716 -480 282828 240 0 FreeSans 448 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 285572 -480 285684 240 0 FreeSans 448 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 288428 -480 288540 240 0 FreeSans 448 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 125636 -480 125748 240 0 FreeSans 448 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 128492 -480 128604 240 0 FreeSans 448 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 131348 -480 131460 240 0 FreeSans 448 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 134204 -480 134316 240 0 FreeSans 448 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 289380 -480 289492 240 0 FreeSans 448 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 290332 -480 290444 240 0 FreeSans 448 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 291284 -480 291396 240 0 FreeSans 448 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 292236 -480 292348 240 0 FreeSans 448 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -478 -342 -168 298654 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -478 -342 298510 -32 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -478 298344 298510 298654 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 298200 -342 298510 298654 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 2709 -822 3019 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 18069 -822 18379 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 33429 -822 33739 74345 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 33429 90103 33739 170745 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 33429 268935 33739 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 48789 -822 49099 74345 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 48789 90103 49099 170745 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 48789 268935 49099 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 64149 -822 64459 74345 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 64149 90103 64459 170745 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 64149 268935 64459 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 79509 -822 79819 170745 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 79509 268935 79819 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 94869 -822 95179 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 110229 -822 110539 97761 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 110229 268935 110539 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 125589 -822 125899 131025 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 125589 268935 125899 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 140949 -822 141259 131025 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 140949 268935 141259 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 156309 -822 156619 131025 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 156309 268935 156619 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 171669 -822 171979 6401 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 171669 158767 171979 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 187029 -822 187339 6401 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 187029 158767 187339 174889 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 187029 191711 187339 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 202389 -822 202699 6401 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 202389 158767 202699 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 217749 -822 218059 6401 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 217749 125367 218059 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 233109 -822 233419 6401 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 233109 125367 233419 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 248469 -822 248779 6401 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 248469 125367 248779 172089 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 248469 187679 248779 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 263829 -822 264139 6401 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 263829 125367 264139 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 279189 -822 279499 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 294549 -822 294859 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 1913 298990 2223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 10913 298990 11223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 19913 298990 20223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 28913 298990 29223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 37913 298990 38223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 46913 298990 47223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 55913 298990 56223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 64913 298990 65223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 73913 298990 74223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 82913 298990 83223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 91913 298990 92223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 100913 298990 101223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 109913 298990 110223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 118913 298990 119223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 127913 298990 128223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 136913 298990 137223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 145913 298990 146223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 154913 298990 155223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 163913 298990 164223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 172913 298990 173223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 181913 298990 182223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 190913 298990 191223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 199913 298990 200223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 208913 298990 209223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 217913 298990 218223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 226913 298990 227223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 235913 298990 236223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 244913 298990 245223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 253913 298990 254223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 262913 298990 263223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 271913 298990 272223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 280913 298990 281223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 289913 298990 290223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -958 -822 -648 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 -822 298990 -512 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 298824 298990 299134 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 298680 -822 298990 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 4569 -822 4879 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 19929 -822 20239 170745 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 19929 268935 20239 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 35289 -822 35599 74345 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 35289 90103 35599 170745 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 35289 268935 35599 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 50649 -822 50959 74345 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 50649 90103 50959 170745 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 50649 268935 50959 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 66009 -822 66319 74345 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 66009 90103 66319 170745 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 66009 268935 66319 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 81369 -822 81679 170745 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 81369 268935 81679 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 96729 -822 97039 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 112089 -822 112399 97761 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 112089 121415 112399 131025 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 112089 268935 112399 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 127449 -822 127759 131025 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 127449 268935 127759 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 142809 -822 143119 131025 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 142809 268935 143119 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 158169 -822 158479 131025 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 158169 268935 158479 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 173529 -822 173839 6401 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 173529 125367 173839 131025 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 173529 158767 173839 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 188889 -822 189199 6401 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 188889 125367 189199 131025 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 188889 191711 189199 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 204249 -822 204559 6401 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 204249 125367 204559 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 219609 -822 219919 6401 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 219609 125367 219919 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 234969 -822 235279 6401 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 234969 125367 235279 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 250329 -822 250639 6401 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 250329 125367 250639 172089 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 250329 187679 250639 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 265689 -822 265999 6401 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 265689 125367 265999 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 281049 -822 281359 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 296409 -822 296719 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 4913 298990 5223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 13913 298990 14223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 22913 298990 23223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 31913 298990 32223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 40913 298990 41223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 49913 298990 50223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 58913 298990 59223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 67913 298990 68223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 76913 298990 77223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 85913 298990 86223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 94913 298990 95223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 103913 298990 104223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 112913 298990 113223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 121913 298990 122223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 130913 298990 131223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 139913 298990 140223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 148913 298990 149223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 157913 298990 158223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 166913 298990 167223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 175913 298990 176223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 184913 298990 185223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 193913 298990 194223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 202913 298990 203223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 211913 298990 212223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 220913 298990 221223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 229913 298990 230223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 238913 298990 239223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 247913 298990 248223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 256913 298990 257223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 265913 298990 266223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 274913 298990 275223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 283913 298990 284223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 292913 298990 293223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 5684 -480 5796 240 0 FreeSans 448 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 6636 -480 6748 240 0 FreeSans 448 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 7588 -480 7700 240 0 FreeSans 448 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 11396 -480 11508 240 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 43764 -480 43876 240 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 46620 -480 46732 240 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 49476 -480 49588 240 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 52332 -480 52444 240 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 55188 -480 55300 240 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 58044 -480 58156 240 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 60900 -480 61012 240 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 63756 -480 63868 240 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 66612 -480 66724 240 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 69468 -480 69580 240 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 15204 -480 15316 240 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 72324 -480 72436 240 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 75180 -480 75292 240 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 78036 -480 78148 240 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 80892 -480 81004 240 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 83748 -480 83860 240 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 86604 -480 86716 240 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 89460 -480 89572 240 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 92316 -480 92428 240 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 95172 -480 95284 240 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 98028 -480 98140 240 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 19012 -480 19124 240 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 100884 -480 100996 240 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 103740 -480 103852 240 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 22820 -480 22932 240 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 26628 -480 26740 240 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 29484 -480 29596 240 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 32340 -480 32452 240 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 35196 -480 35308 240 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 38052 -480 38164 240 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 40908 -480 41020 240 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 8540 -480 8652 240 0 FreeSans 448 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 12348 -480 12460 240 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 44716 -480 44828 240 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 47572 -480 47684 240 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 50428 -480 50540 240 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 53284 -480 53396 240 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 56140 -480 56252 240 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 58996 -480 59108 240 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 61852 -480 61964 240 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 64708 -480 64820 240 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 67564 -480 67676 240 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 70420 -480 70532 240 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 16156 -480 16268 240 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 73276 -480 73388 240 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 76132 -480 76244 240 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 78988 -480 79100 240 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 81844 -480 81956 240 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 84700 -480 84812 240 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 87556 -480 87668 240 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 90412 -480 90524 240 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 93268 -480 93380 240 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 96124 -480 96236 240 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 98980 -480 99092 240 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 19964 -480 20076 240 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 101836 -480 101948 240 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 104692 -480 104804 240 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 23772 -480 23884 240 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 27580 -480 27692 240 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 30436 -480 30548 240 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 33292 -480 33404 240 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 36148 -480 36260 240 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 39004 -480 39116 240 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 41860 -480 41972 240 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 13300 -480 13412 240 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 45668 -480 45780 240 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 48524 -480 48636 240 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 51380 -480 51492 240 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 54236 -480 54348 240 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 57092 -480 57204 240 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 59948 -480 60060 240 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 62804 -480 62916 240 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 65660 -480 65772 240 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 68516 -480 68628 240 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 71372 -480 71484 240 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 17108 -480 17220 240 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 74228 -480 74340 240 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 77084 -480 77196 240 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 79940 -480 80052 240 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 82796 -480 82908 240 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 85652 -480 85764 240 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 88508 -480 88620 240 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 91364 -480 91476 240 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 94220 -480 94332 240 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 97076 -480 97188 240 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 99932 -480 100044 240 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 20916 -480 21028 240 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 102788 -480 102900 240 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 105644 -480 105756 240 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 24724 -480 24836 240 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 28532 -480 28644 240 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 31388 -480 31500 240 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 34244 -480 34356 240 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 37100 -480 37212 240 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 39956 -480 40068 240 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 42812 -480 42924 240 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 14252 -480 14364 240 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 18060 -480 18172 240 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 21868 -480 21980 240 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 25676 -480 25788 240 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 9492 -480 9604 240 0 FreeSans 448 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 10444 -480 10556 240 0 FreeSans 448 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 93135 101161 93135 101161 0 vdd
rlabel via4 85455 95161 85455 95161 0 vss
rlabel metal2 163156 126959 163156 126959 0 diego_clk
rlabel metal2 225260 128793 225260 128793 0 diego_io_in_all38\[10\]
rlabel metal2 225932 128429 225932 128429 0 diego_io_in_all38\[11\]
rlabel metal2 226604 128765 226604 128765 0 diego_io_in_all38\[12\]
rlabel metal2 227276 128737 227276 128737 0 diego_io_in_all38\[13\]
rlabel metal2 247156 126175 247156 126175 0 diego_io_in_all38\[14\]
rlabel metal2 248276 126147 248276 126147 0 diego_io_in_all38\[15\]
rlabel metal2 229292 128653 229292 128653 0 diego_io_in_all38\[16\]
rlabel metal2 229964 129185 229964 129185 0 diego_io_in_all38\[17\]
rlabel metal3 247884 128352 247884 128352 0 diego_io_in_all38\[18\]
rlabel metal3 247940 128268 247940 128268 0 diego_io_in_all38\[19\]
rlabel metal2 231980 129101 231980 129101 0 diego_io_in_all38\[20\]
rlabel metal2 232652 129521 232652 129521 0 diego_io_in_all38\[21\]
rlabel metal2 233324 129661 233324 129661 0 diego_io_in_all38\[22\]
rlabel metal2 233996 129633 233996 129633 0 diego_io_in_all38\[23\]
rlabel metal2 234668 129577 234668 129577 0 diego_io_in_all38\[24\]
rlabel metal2 235340 129073 235340 129073 0 diego_io_in_all38\[25\]
rlabel metal2 236012 129549 236012 129549 0 diego_io_in_all38\[26\]
rlabel metal2 236684 129689 236684 129689 0 diego_io_in_all38\[27\]
rlabel metal2 237356 129493 237356 129493 0 diego_io_in_all38\[28\]
rlabel metal2 238028 128401 238028 128401 0 diego_io_in_all38\[29\]
rlabel metal2 238700 128373 238700 128373 0 diego_io_in_all38\[30\]
rlabel metal2 239372 128345 239372 128345 0 diego_io_in_all38\[31\]
rlabel metal2 240044 129521 240044 129521 0 diego_io_in_all38\[32\]
rlabel metal2 240716 128317 240716 128317 0 diego_io_in_all38\[33\]
rlabel metal2 269556 126623 269556 126623 0 diego_io_in_all38\[34\]
rlabel metal2 270676 125755 270676 125755 0 diego_io_in_all38\[35\]
rlabel metal2 271796 125727 271796 125727 0 diego_io_in_all38\[36\]
rlabel metal2 272916 125699 272916 125699 0 diego_io_in_all38\[37\]
rlabel metal2 222572 129577 222572 129577 0 diego_io_in_all38\[6\]
rlabel metal2 223244 129633 223244 129633 0 diego_io_in_all38\[7\]
rlabel metal2 223916 129297 223916 129297 0 diego_io_in_all38\[8\]
rlabel metal2 224588 129605 224588 129605 0 diego_io_in_all38\[9\]
rlabel metal2 202356 126959 202356 126959 0 diego_io_oeb\[0\]
rlabel metal2 203756 129577 203756 129577 0 diego_io_oeb\[10\]
rlabel metal2 214676 126959 214676 126959 0 diego_io_oeb\[11\]
rlabel metal2 215796 125727 215796 125727 0 diego_io_oeb\[12\]
rlabel metal2 205772 128233 205772 128233 0 diego_io_oeb\[13\]
rlabel metal2 206444 128205 206444 128205 0 diego_io_oeb\[14\]
rlabel metal2 207116 128429 207116 128429 0 diego_io_oeb\[15\]
rlabel metal2 207788 128765 207788 128765 0 diego_io_oeb\[16\]
rlabel metal2 208460 128737 208460 128737 0 diego_io_oeb\[17\]
rlabel metal2 222516 126175 222516 126175 0 diego_io_oeb\[18\]
rlabel metal2 223636 126147 223636 126147 0 diego_io_oeb\[19\]
rlabel metal2 203476 126567 203476 126567 0 diego_io_oeb\[1\]
rlabel metal2 210476 129549 210476 129549 0 diego_io_oeb\[20\]
rlabel metal2 211148 128653 211148 128653 0 diego_io_oeb\[21\]
rlabel metal2 211820 129521 211820 129521 0 diego_io_oeb\[22\]
rlabel metal2 212492 129073 212492 129073 0 diego_io_oeb\[23\]
rlabel metal2 213164 128401 213164 128401 0 diego_io_oeb\[24\]
rlabel metal2 213836 128373 213836 128373 0 diego_io_oeb\[25\]
rlabel metal2 214508 128345 214508 128345 0 diego_io_oeb\[26\]
rlabel metal2 215180 128317 215180 128317 0 diego_io_oeb\[27\]
rlabel metal2 215852 128289 215852 128289 0 diego_io_oeb\[28\]
rlabel metal2 234836 125727 234836 125727 0 diego_io_oeb\[29\]
rlabel metal2 198380 129073 198380 129073 0 diego_io_oeb\[2\]
rlabel metal2 235956 125699 235956 125699 0 diego_io_oeb\[30\]
rlabel metal2 237076 125587 237076 125587 0 diego_io_oeb\[31\]
rlabel metal2 199052 128373 199052 128373 0 diego_io_oeb\[3\]
rlabel metal2 199724 128681 199724 128681 0 diego_io_oeb\[4\]
rlabel metal2 200396 128345 200396 128345 0 diego_io_oeb\[5\]
rlabel metal2 201068 128317 201068 128317 0 diego_io_oeb\[6\]
rlabel metal2 201740 128653 201740 128653 0 diego_io_oeb\[7\]
rlabel metal2 202412 128289 202412 128289 0 diego_io_oeb\[8\]
rlabel metal2 203084 128793 203084 128793 0 diego_io_oeb\[9\]
rlabel metal2 166516 125699 166516 125699 0 diego_io_out\[0\]
rlabel metal2 177716 126763 177716 126763 0 diego_io_out\[10\]
rlabel metal2 178836 127015 178836 127015 0 diego_io_out\[11\]
rlabel metal2 179956 127043 179956 127043 0 diego_io_out\[12\]
rlabel metal3 182672 128884 182672 128884 0 diego_io_out\[13\]
rlabel metal3 183568 128940 183568 128940 0 diego_io_out\[14\]
rlabel metal3 184464 128828 184464 128828 0 diego_io_out\[15\]
rlabel metal3 185360 128884 185360 128884 0 diego_io_out\[16\]
rlabel metal2 186956 129297 186956 129297 0 diego_io_out\[17\]
rlabel metal2 186676 125923 186676 125923 0 diego_io_out\[18\]
rlabel metal2 188300 128863 188300 128863 0 diego_io_out\[19\]
rlabel metal2 167636 125727 167636 125727 0 diego_io_out\[1\]
rlabel metal2 188937 130060 188937 130060 0 diego_io_out\[20\]
rlabel metal2 189840 128884 189840 128884 0 diego_io_out\[21\]
rlabel metal3 190736 128884 190736 128884 0 diego_io_out\[22\]
rlabel metal3 191632 128828 191632 128828 0 diego_io_out\[23\]
rlabel metal2 191660 128429 191660 128429 0 diego_io_out\[24\]
rlabel metal2 192332 128233 192332 128233 0 diego_io_out\[25\]
rlabel metal2 195636 125615 195636 125615 0 diego_io_out\[26\]
rlabel metal2 196756 125587 196756 125587 0 diego_io_out\[27\]
rlabel metal2 197876 125559 197876 125559 0 diego_io_out\[28\]
rlabel metal2 198996 125867 198996 125867 0 diego_io_out\[29\]
rlabel metal2 168756 125755 168756 125755 0 diego_io_out\[2\]
rlabel metal2 200116 127015 200116 127015 0 diego_io_out\[30\]
rlabel metal2 201236 126987 201236 126987 0 diego_io_out\[31\]
rlabel metal2 177548 129521 177548 129521 0 diego_io_out\[3\]
rlabel metal2 178220 129549 178220 129549 0 diego_io_out\[4\]
rlabel metal2 178892 129577 178892 129577 0 diego_io_out\[5\]
rlabel metal2 179564 128317 179564 128317 0 diego_io_out\[6\]
rlabel metal2 180236 129493 180236 129493 0 diego_io_out\[7\]
rlabel metal2 175476 126539 175476 126539 0 diego_io_out\[8\]
rlabel metal2 176596 125895 176596 125895 0 diego_io_out\[9\]
rlabel metal3 286881 3556 286881 3556 0 io_in[0]
rlabel metal3 296653 201796 296653 201796 0 io_in[10]
rlabel metal3 296625 221620 296625 221620 0 io_in[11]
rlabel metal3 296597 241444 296597 241444 0 io_in[12]
rlabel metal3 296569 261268 296569 261268 0 io_in[13]
rlabel metal3 296541 281092 296541 281092 0 io_in[14]
rlabel metal2 292348 227969 292348 227969 0 io_in[15]
rlabel metal2 259252 296541 259252 296541 0 io_in[16]
rlabel metal3 225428 295092 225428 295092 0 io_in[17]
rlabel metal2 222236 160867 222236 160867 0 io_in[18]
rlabel metal2 93884 227619 93884 227619 0 io_in[19]
rlabel metal3 286965 23380 286965 23380 0 io_in[1]
rlabel metal2 93660 228760 93660 228760 0 io_in[20]
rlabel metal2 93772 229929 93772 229929 0 io_in[21]
rlabel metal2 60788 296597 60788 296597 0 io_in[22]
rlabel metal2 27580 296541 27580 296541 0 io_in[23]
rlabel metal3 1995 293580 1995 293580 0 io_in[24]
rlabel metal3 1659 272412 1659 272412 0 io_in[25]
rlabel metal3 2023 251244 2023 251244 0 io_in[26]
rlabel metal3 2051 230076 2051 230076 0 io_in[27]
rlabel metal3 2079 208908 2079 208908 0 io_in[28]
rlabel metal3 2583 187740 2583 187740 0 io_in[29]
rlabel metal3 273007 140644 273007 140644 0 io_in[2]
rlabel metal3 2107 166572 2107 166572 0 io_in[30]
rlabel metal3 1351 145404 1351 145404 0 io_in[31]
rlabel metal3 29113 142660 29113 142660 0 io_in[32]
rlabel metal3 1687 103180 1687 103180 0 io_in[33]
rlabel metal3 2079 82012 2079 82012 0 io_in[34]
rlabel metal3 2051 60844 2051 60844 0 io_in[35]
rlabel metal3 1659 39676 1659 39676 0 io_in[36]
rlabel metal3 1995 18452 1995 18452 0 io_in[37]
rlabel metal3 273063 141988 273063 141988 0 io_in[3]
rlabel metal3 273427 143332 273427 143332 0 io_in[4]
rlabel metal3 273455 144676 273455 144676 0 io_in[5]
rlabel metal3 273483 146020 273483 146020 0 io_in[6]
rlabel metal3 270935 147364 270935 147364 0 io_in[7]
rlabel metal3 271383 148708 271383 148708 0 io_in[8]
rlabel metal3 271355 150052 271355 150052 0 io_in[9]
rlabel metal3 272979 138852 272979 138852 0 io_oeb[0]
rlabel metal3 271327 152292 271327 152292 0 io_oeb[10]
rlabel metal3 271691 153636 271691 153636 0 io_oeb[11]
rlabel metal3 271271 154980 271271 154980 0 io_oeb[12]
rlabel metal3 272531 156324 272531 156324 0 io_oeb[13]
rlabel metal3 286881 294308 286881 294308 0 io_oeb[14]
rlabel metal2 269976 297836 269976 297836 0 io_oeb[15]
rlabel metal2 237188 296597 237188 296597 0 io_oeb[16]
rlabel metal2 222908 160839 222908 160839 0 io_oeb[17]
rlabel metal2 171108 296541 171108 296541 0 io_oeb[18]
rlabel metal2 92540 160643 92540 160643 0 io_oeb[19]
rlabel metal3 273371 140196 273371 140196 0 io_oeb[1]
rlabel metal2 104804 296681 104804 296681 0 io_oeb[20]
rlabel metal2 71820 296625 71820 296625 0 io_oeb[21]
rlabel metal2 38724 296541 38724 296541 0 io_oeb[22]
rlabel metal3 17773 156660 17773 156660 0 io_oeb[23]
rlabel metal3 17745 154980 17745 154980 0 io_oeb[24]
rlabel metal3 2863 258300 2863 258300 0 io_oeb[25]
rlabel metal3 2891 237132 2891 237132 0 io_oeb[26]
rlabel metal3 2919 215964 2919 215964 0 io_oeb[27]
rlabel metal3 3283 194796 3283 194796 0 io_oeb[28]
rlabel metal3 1687 173628 1687 173628 0 io_oeb[29]
rlabel metal3 273399 141540 273399 141540 0 io_oeb[2]
rlabel metal3 1155 152460 1155 152460 0 io_oeb[30]
rlabel metal3 14231 131292 14231 131292 0 io_oeb[31]
rlabel metal3 29085 141540 29085 141540 0 io_oeb[32]
rlabel metal3 2107 89012 2107 89012 0 io_oeb[33]
rlabel metal3 1267 67900 1267 67900 0 io_oeb[34]
rlabel metal3 1211 46732 1211 46732 0 io_oeb[35]
rlabel metal3 2835 25564 2835 25564 0 io_oeb[36]
rlabel metal3 1155 4396 1155 4396 0 io_oeb[37]
rlabel metal3 270963 142884 270963 142884 0 io_oeb[3]
rlabel metal3 270907 144228 270907 144228 0 io_oeb[4]
rlabel metal3 296653 116004 296653 116004 0 io_oeb[5]
rlabel metal3 270879 146916 270879 146916 0 io_oeb[6]
rlabel metal3 270851 148260 270851 148260 0 io_oeb[7]
rlabel metal3 270935 149604 270935 149604 0 io_oeb[8]
rlabel metal3 273371 150948 273371 150948 0 io_oeb[9]
rlabel metal3 270879 151844 270879 151844 0 io_out[10]
rlabel metal3 273791 153188 273791 153188 0 io_out[11]
rlabel metal3 271299 154532 271299 154532 0 io_out[12]
rlabel metal3 274211 155876 274211 155876 0 io_out[13]
rlabel metal3 270851 157220 270851 157220 0 io_out[14]
rlabel metal2 281316 296541 281316 296541 0 io_out[15]
rlabel metal2 248220 296569 248220 296569 0 io_out[16]
rlabel metal2 215124 232281 215124 232281 0 io_out[17]
rlabel metal2 182140 296569 182140 296569 0 io_out[18]
rlabel metal2 93212 160867 93212 160867 0 io_out[19]
rlabel metal2 115836 296653 115836 296653 0 io_out[20]
rlabel metal2 82852 296737 82852 296737 0 io_out[21]
rlabel metal2 49756 296569 49756 296569 0 io_out[22]
rlabel metal2 16548 227521 16548 227521 0 io_out[23]
rlabel metal3 1155 286524 1155 286524 0 io_out[24]
rlabel metal3 1183 265356 1183 265356 0 io_out[25]
rlabel metal3 1211 244188 1211 244188 0 io_out[26]
rlabel metal3 1239 223020 1239 223020 0 io_out[27]
rlabel metal3 3255 201852 3255 201852 0 io_out[28]
rlabel metal3 1267 180684 1267 180684 0 io_out[29]
rlabel metal3 3311 159516 3311 159516 0 io_out[30]
rlabel metal3 1155 138460 1155 138460 0 io_out[31]
rlabel metal3 1295 117292 1295 117292 0 io_out[32]
rlabel metal3 3255 96012 3255 96012 0 io_out[33]
rlabel metal3 3675 74844 3675 74844 0 io_out[34]
rlabel metal3 1239 53732 1239 53732 0 io_out[35]
rlabel metal3 2023 32620 2023 32620 0 io_out[36]
rlabel metal3 1183 11452 1183 11452 0 io_out[37]
rlabel metal3 270963 149156 270963 149156 0 io_out[8]
rlabel metal3 270907 150500 270907 150500 0 io_out[9]
rlabel metal2 143948 66101 143948 66101 0 la_data_in[10]
rlabel metal2 144620 129521 144620 129521 0 la_data_in[11]
rlabel metal2 140980 1127 140980 1127 0 la_data_in[12]
rlabel metal2 143836 1351 143836 1351 0 la_data_in[13]
rlabel metal2 146601 130060 146601 130060 0 la_data_in[14]
rlabel metal3 148372 2100 148372 2100 0 la_data_in[15]
rlabel metal2 152292 1323 152292 1323 0 la_data_in[16]
rlabel metal2 155148 64603 155148 64603 0 la_data_in[17]
rlabel metal2 158004 1575 158004 1575 0 la_data_in[18]
rlabel metal2 149996 129493 149996 129493 0 la_data_in[19]
rlabel metal2 163716 1239 163716 1239 0 la_data_in[20]
rlabel metal2 166572 1211 166572 1211 0 la_data_in[21]
rlabel metal2 152012 66101 152012 66101 0 la_data_in[22]
rlabel metal2 152684 66073 152684 66073 0 la_data_in[23]
rlabel metal3 274127 130788 274127 130788 0 la_data_in[48]
rlabel metal2 246652 1995 246652 1995 0 la_data_in[49]
rlabel metal2 249396 3283 249396 3283 0 la_data_in[50]
rlabel metal3 274015 132132 274015 132132 0 la_data_in[51]
rlabel metal2 255220 2023 255220 2023 0 la_data_in[52]
rlabel metal2 258076 1575 258076 1575 0 la_data_in[53]
rlabel metal2 260820 3311 260820 3311 0 la_data_in[54]
rlabel metal2 263732 1603 263732 1603 0 la_data_in[55]
rlabel metal2 266644 1631 266644 1631 0 la_data_in[56]
rlabel metal2 269388 3675 269388 3675 0 la_data_in[57]
rlabel metal2 272356 1155 272356 1155 0 la_data_in[58]
rlabel metal3 269948 135681 269948 135681 0 la_data_in[59]
rlabel metal3 273959 136164 273959 136164 0 la_data_in[60]
rlabel metal2 280812 1351 280812 1351 0 la_data_in[61]
rlabel metal2 283668 1183 283668 1183 0 la_data_in[62]
rlabel metal2 286524 1155 286524 1155 0 la_data_in[63]
rlabel metal2 129556 1155 129556 1155 0 la_data_in[8]
rlabel metal2 143276 129493 143276 129493 0 la_data_in[9]
rlabel metal2 70700 129493 70700 129493 0 pawel_io_in_all38\[25\]
rlabel metal2 24444 106043 24444 106043 0 pawel_io_in_all38\[26\]
rlabel metal2 72044 129521 72044 129521 0 pawel_io_in_all38\[27\]
rlabel metal2 35868 106071 35868 106071 0 pawel_io_in_all38\[28\]
rlabel metal2 73388 118629 73388 118629 0 pawel_io_in_all38\[29\]
rlabel metal2 47292 106127 47292 106127 0 pawel_io_in_all38\[30\]
rlabel metal2 74732 118685 74732 118685 0 pawel_io_in_all38\[31\]
rlabel metal2 58716 106211 58716 106211 0 pawel_io_in_all38\[32\]
rlabel metal2 64428 105819 64428 105819 0 pawel_io_in_all38\[33\]
rlabel metal2 70140 117019 70140 117019 0 pawel_io_in_all38\[34\]
rlabel metal3 76636 128884 76636 128884 0 pawel_io_in_all38\[35\]
rlabel metal2 81564 105819 81564 105819 0 pawel_io_in_all38\[36\]
rlabel metal2 87276 105763 87276 105763 0 pawel_io_in_all38\[37\]
rlabel metal2 37100 118153 37100 118153 0 pawel_io_oeb\[0\]
rlabel metal2 57260 118713 57260 118713 0 pawel_io_oeb\[10\]
rlabel metal2 83468 105679 83468 105679 0 pawel_io_oeb\[11\]
rlabel metal2 61292 118153 61292 118153 0 pawel_io_oeb\[12\]
rlabel metal2 26348 105707 26348 105707 0 pawel_io_oeb\[1\]
rlabel metal2 32060 105763 32060 105763 0 pawel_io_oeb\[2\]
rlabel metal2 37772 105623 37772 105623 0 pawel_io_oeb\[3\]
rlabel metal2 43484 105819 43484 105819 0 pawel_io_oeb\[4\]
rlabel metal2 49196 105819 49196 105819 0 pawel_io_oeb\[5\]
rlabel metal3 49588 128884 49588 128884 0 pawel_io_oeb\[6\]
rlabel metal2 51212 129297 51212 129297 0 pawel_io_oeb\[7\]
rlabel metal2 66332 105707 66332 105707 0 pawel_io_oeb\[8\]
rlabel metal2 72044 105763 72044 105763 0 pawel_io_oeb\[9\]
rlabel metal2 22540 105679 22540 105679 0 pawel_io_out\[0\]
rlabel metal2 57932 118265 57932 118265 0 pawel_io_out\[10\]
rlabel metal2 85372 105651 85372 105651 0 pawel_io_out\[11\]
rlabel metal2 61964 129633 61964 129633 0 pawel_io_out\[12\]
rlabel metal2 28252 105735 28252 105735 0 pawel_io_out\[1\]
rlabel metal2 33964 117019 33964 117019 0 pawel_io_out\[2\]
rlabel metal2 39676 105791 39676 105791 0 pawel_io_out\[3\]
rlabel metal2 45605 130060 45605 130060 0 pawel_io_out\[4\]
rlabel metal2 51100 105791 51100 105791 0 pawel_io_out\[5\]
rlabel metal2 49868 118181 49868 118181 0 pawel_io_out\[6\]
rlabel metal2 62524 105791 62524 105791 0 pawel_io_out\[7\]
rlabel metal2 53900 129549 53900 129549 0 pawel_io_out\[8\]
rlabel metal2 73948 105791 73948 105791 0 pawel_io_out\[9\]
rlabel metal2 35084 129521 35084 129521 0 pawel_mux_rst
rlabel metal2 235900 167965 235900 167965 0 solos_clk
rlabel metal2 237244 167993 237244 167993 0 solos_gpio_ready
rlabel metal2 259868 162519 259868 162519 0 solos_io_in_all38\[10\]
rlabel metal2 259196 161287 259196 161287 0 solos_io_in_all38\[11\]
rlabel metal2 258524 161259 258524 161259 0 solos_io_in_all38\[12\]
rlabel metal2 257852 162967 257852 162967 0 solos_io_in_all38\[13\]
rlabel metal2 250684 166705 250684 166705 0 solos_io_in_all38\[14\]
rlabel metal2 250012 167153 250012 167153 0 solos_io_in_all38\[15\]
rlabel metal2 249340 166733 249340 166733 0 solos_io_in_all38\[16\]
rlabel metal2 248668 167965 248668 167965 0 solos_io_in_all38\[17\]
rlabel metal2 247996 168021 247996 168021 0 solos_io_in_all38\[18\]
rlabel metal2 247324 167181 247324 167181 0 solos_io_in_all38\[19\]
rlabel metal2 246652 167125 246652 167125 0 solos_io_in_all38\[20\]
rlabel metal2 261212 164199 261212 164199 0 solos_io_in_all38\[8\]
rlabel metal2 260540 161735 260540 161735 0 solos_io_in_all38\[9\]
rlabel metal2 245980 168945 245980 168945 0 solos_io_out\[0\]
rlabel metal3 236796 165788 236796 165788 0 solos_io_out\[10\]
rlabel metal3 236124 165844 236124 165844 0 solos_io_out\[11\]
rlabel metal2 237916 168133 237916 168133 0 solos_io_out\[12\]
rlabel metal2 245308 168973 245308 168973 0 solos_io_out\[1\]
rlabel metal3 242172 167188 242172 167188 0 solos_io_out\[2\]
rlabel metal2 239036 163975 239036 163975 0 solos_io_out\[3\]
rlabel metal2 238364 163835 238364 163835 0 solos_io_out\[4\]
rlabel metal2 237692 163779 237692 163779 0 solos_io_out\[5\]
rlabel metal2 237020 163807 237020 163807 0 solos_io_out\[6\]
rlabel metal2 236348 163863 236348 163863 0 solos_io_out\[7\]
rlabel metal2 235676 163135 235676 163135 0 solos_io_out\[8\]
rlabel metal2 235004 163079 235004 163079 0 solos_io_out\[9\]
rlabel metal2 236572 165865 236572 165865 0 solos_rst
rlabel metal3 102452 167188 102452 167188 0 trzf2_clk
rlabel metal2 163436 166285 163436 166285 0 trzf2_io_in\[18\]
rlabel metal2 134204 161287 134204 161287 0 trzf2_io_in\[19\]
rlabel metal2 133532 161315 133532 161315 0 trzf2_io_in\[20\]
rlabel metal2 132860 161343 132860 161343 0 trzf2_io_in\[21\]
rlabel metal2 132188 161371 132188 161371 0 trzf2_io_in\[22\]
rlabel metal2 131516 161399 131516 161399 0 trzf2_io_in\[23\]
rlabel metal2 130844 161427 130844 161427 0 trzf2_io_in\[24\]
rlabel metal2 130172 161063 130172 161063 0 trzf2_io_in\[25\]
rlabel metal2 129500 160839 129500 160839 0 trzf2_io_in\[26\]
rlabel metal2 128828 161287 128828 161287 0 trzf2_io_in\[27\]
rlabel metal2 128156 160867 128156 160867 0 trzf2_io_in\[28\]
rlabel metal2 132300 165592 132300 165592 0 trzf2_io_in\[29\]
rlabel metal2 126812 160895 126812 160895 0 trzf2_io_in\[30\]
rlabel metal2 131628 165564 131628 165564 0 trzf2_io_in\[31\]
rlabel metal2 144620 165949 144620 165949 0 trzf2_io_in\[32\]
rlabel metal2 129948 165144 129948 165144 0 trzf2_io_in\[33\]
rlabel metal2 141932 166005 141932 166005 0 trzf2_io_in\[34\]
rlabel metal3 106484 163772 106484 163772 0 trzf2_la_in\[10\]
rlabel metal2 106988 166733 106988 166733 0 trzf2_la_in\[11\]
rlabel metal2 105644 168693 105644 168693 0 trzf2_la_in\[12\]
rlabel metal3 118608 163772 118608 163772 0 trzf2_la_in\[1\]
rlabel metal2 110012 163807 110012 163807 0 trzf2_la_in\[2\]
rlabel metal2 109340 163835 109340 163835 0 trzf2_la_in\[3\]
rlabel metal2 108668 163863 108668 163863 0 trzf2_la_in\[4\]
rlabel metal2 107996 163891 107996 163891 0 trzf2_la_in\[5\]
rlabel metal2 107324 163919 107324 163919 0 trzf2_la_in\[6\]
rlabel metal2 106652 163947 106652 163947 0 trzf2_la_in\[7\]
rlabel metal2 105980 163667 105980 163667 0 trzf2_la_in\[8\]
rlabel metal3 107492 168028 107492 168028 0 trzf2_la_in\[9\]
rlabel metal2 113372 160895 113372 160895 0 trzf2_o_gpout\[0\]
rlabel metal2 112700 161259 112700 161259 0 trzf2_o_gpout\[1\]
rlabel metal2 121772 168805 121772 168805 0 trzf2_o_gpout\[2\]
rlabel metal2 121436 161679 121436 161679 0 trzf2_o_hsync
rlabel metal2 120092 161707 120092 161707 0 trzf2_o_rgb\[0\]
rlabel metal2 119420 161007 119420 161007 0 trzf2_o_rgb\[1\]
rlabel metal2 118748 161035 118748 161035 0 trzf2_o_rgb\[2\]
rlabel metal2 118076 164199 118076 164199 0 trzf2_o_rgb\[3\]
rlabel metal2 117404 164227 117404 164227 0 trzf2_o_rgb\[4\]
rlabel metal2 116732 164255 116732 164255 0 trzf2_o_rgb\[5\]
rlabel metal2 116060 164283 116060 164283 0 trzf2_o_tex_csb
rlabel metal2 114044 160867 114044 160867 0 trzf2_o_tex_oeb0
rlabel metal3 120932 168644 120932 168644 0 trzf2_o_tex_out0
rlabel metal2 128492 165865 128492 165865 0 trzf2_o_tex_sclk
rlabel metal2 120764 160951 120764 160951 0 trzf2_o_vsync
rlabel metal2 104300 168665 104300 168665 0 trzf2_rst
rlabel metal2 22932 169225 22932 169225 0 trzf_clk
rlabel metal2 83412 165865 83412 165865 0 trzf_io_in\[18\]
rlabel metal2 82068 165893 82068 165893 0 trzf_io_in\[19\]
rlabel metal2 70980 163520 70980 163520 0 trzf_io_in\[20\]
rlabel metal2 64988 160895 64988 160895 0 trzf_io_in\[21\]
rlabel metal2 64316 160923 64316 160923 0 trzf_io_in\[22\]
rlabel metal2 63644 160951 63644 160951 0 trzf_io_in\[23\]
rlabel metal2 62972 161007 62972 161007 0 trzf_io_in\[24\]
rlabel metal2 62300 161035 62300 161035 0 trzf_io_in\[25\]
rlabel metal2 61628 164199 61628 164199 0 trzf_io_in\[26\]
rlabel metal2 60956 164283 60956 164283 0 trzf_io_in\[27\]
rlabel metal2 60284 164311 60284 164311 0 trzf_io_in\[28\]
rlabel metal2 59612 163359 59612 163359 0 trzf_io_in\[29\]
rlabel metal2 58940 163387 58940 163387 0 trzf_io_in\[30\]
rlabel metal2 58268 163415 58268 163415 0 trzf_io_in\[31\]
rlabel metal2 57596 163471 57596 163471 0 trzf_io_in\[32\]
rlabel metal3 60088 167020 60088 167020 0 trzf_io_in\[33\]
rlabel metal2 61908 165865 61908 165865 0 trzf_io_in\[34\]
rlabel metal2 36764 160895 36764 160895 0 trzf_la_in\[10\]
rlabel metal2 26964 168385 26964 168385 0 trzf_la_in\[11\]
rlabel metal2 25620 165893 25620 165893 0 trzf_la_in\[12\]
rlabel metal2 42812 160643 42812 160643 0 trzf_la_in\[1\]
rlabel metal2 39060 165949 39060 165949 0 trzf_la_in\[2\]
rlabel metal2 37716 165921 37716 165921 0 trzf_la_in\[3\]
rlabel metal2 36372 166061 36372 166061 0 trzf_la_in\[4\]
rlabel metal2 35028 165865 35028 165865 0 trzf_la_in\[5\]
rlabel metal2 39452 160643 39452 160643 0 trzf_la_in\[6\]
rlabel metal2 38780 161259 38780 161259 0 trzf_la_in\[7\]
rlabel metal2 38108 162099 38108 162099 0 trzf_la_in\[8\]
rlabel metal2 37436 160923 37436 160923 0 trzf_la_in\[9\]
rlabel metal2 45500 161035 45500 161035 0 trzf_o_gpout\[0\]
rlabel metal2 44828 160643 44828 160643 0 trzf_o_gpout\[1\]
rlabel metal2 44156 161063 44156 161063 0 trzf_o_gpout\[2\]
rlabel metal2 60564 168469 60564 168469 0 trzf_o_hsync
rlabel metal2 57876 168805 57876 168805 0 trzf_o_rgb\[0\]
rlabel metal3 54040 167188 54040 167188 0 trzf_o_rgb\[1\]
rlabel metal2 50876 163835 50876 163835 0 trzf_o_rgb\[2\]
rlabel metal2 50204 163863 50204 163863 0 trzf_o_rgb\[3\]
rlabel metal2 49532 161483 49532 161483 0 trzf_o_rgb\[4\]
rlabel metal3 50008 167188 50008 167188 0 trzf_o_rgb\[5\]
rlabel metal3 49000 167244 49000 167244 0 trzf_o_tex_csb
rlabel metal2 45983 170044 45983 170044 0 trzf_o_tex_oeb0
rlabel metal2 46956 167188 46956 167188 0 trzf_o_tex_out0
rlabel metal3 47992 167188 47992 167188 0 trzf_o_tex_sclk
rlabel metal2 59220 168385 59220 168385 0 trzf_o_vsync
rlabel metal2 24276 165865 24276 165865 0 trzf_rst
rlabel metal2 82796 128653 82796 128653 0 uri_clk
rlabel metal2 84812 128681 84812 128681 0 uri_io_in\[0\]
rlabel metal2 109228 125923 109228 125923 0 uri_io_in\[10\]
rlabel metal2 109900 125559 109900 125559 0 uri_io_in\[11\]
rlabel metal2 109004 128401 109004 128401 0 uri_io_in\[12\]
rlabel metal2 111139 130060 111139 130060 0 uri_io_in\[13\]
rlabel metal2 111916 125923 111916 125923 0 uri_io_in\[14\]
rlabel metal3 113820 128884 113820 128884 0 uri_io_in\[15\]
rlabel metal2 117068 129325 117068 129325 0 uri_io_in\[16\]
rlabel metal2 119049 130060 119049 130060 0 uri_io_in\[17\]
rlabel metal2 121100 129549 121100 129549 0 uri_io_in\[18\]
rlabel metal2 123116 129521 123116 129521 0 uri_io_in\[19\]
rlabel metal2 86828 128709 86828 128709 0 uri_io_in\[1\]
rlabel metal2 115948 126959 115948 126959 0 uri_io_in\[20\]
rlabel metal2 116620 126539 116620 126539 0 uri_io_in\[21\]
rlabel metal2 117292 125699 117292 125699 0 uri_io_in\[22\]
rlabel metal2 117964 125783 117964 125783 0 uri_io_in\[23\]
rlabel metal2 118636 127127 118636 127127 0 uri_io_in\[24\]
rlabel metal2 119308 127071 119308 127071 0 uri_io_in\[25\]
rlabel metal2 119980 125839 119980 125839 0 uri_io_in\[26\]
rlabel metal2 128492 129465 128492 129465 0 uri_io_in\[27\]
rlabel metal2 129164 129633 129164 129633 0 uri_io_in\[28\]
rlabel metal2 129836 129577 129836 129577 0 uri_io_in\[29\]
rlabel metal2 88844 128737 88844 128737 0 uri_io_in\[2\]
rlabel metal2 130508 128345 130508 128345 0 uri_io_in\[30\]
rlabel metal2 131180 128317 131180 128317 0 uri_io_in\[31\]
rlabel metal2 131852 128261 131852 128261 0 uri_io_in\[32\]
rlabel metal2 132524 129689 132524 129689 0 uri_io_in\[33\]
rlabel metal2 133196 128233 133196 128233 0 uri_io_in\[34\]
rlabel metal2 133868 129549 133868 129549 0 uri_io_in\[35\]
rlabel metal2 134540 129661 134540 129661 0 uri_io_in\[36\]
rlabel metal2 135212 129521 135212 129521 0 uri_io_in\[37\]
rlabel metal2 104524 125867 104524 125867 0 uri_io_in\[3\]
rlabel metal2 92876 128765 92876 128765 0 uri_io_in\[4\]
rlabel metal2 94892 128205 94892 128205 0 uri_io_in\[5\]
rlabel metal2 96908 129605 96908 129605 0 uri_io_in\[6\]
rlabel metal2 107212 126679 107212 126679 0 uri_io_in\[7\]
rlabel metal2 107884 127099 107884 127099 0 uri_io_in\[8\]
rlabel metal2 108556 126091 108556 126091 0 uri_io_in\[9\]
rlabel metal2 109452 126539 109452 126539 0 uri_io_oeb\[10\]
rlabel metal2 91532 129633 91532 129633 0 uri_io_oeb\[11\]
rlabel metal2 93548 129101 93548 129101 0 uri_io_oeb\[12\]
rlabel metal2 95564 129661 95564 129661 0 uri_io_oeb\[13\]
rlabel metal2 97580 129689 97580 129689 0 uri_io_oeb\[14\]
rlabel metal2 99596 129129 99596 129129 0 uri_io_oeb\[15\]
rlabel metal2 101612 129157 101612 129157 0 uri_io_oeb\[16\]
rlabel metal2 103628 128317 103628 128317 0 uri_io_oeb\[17\]
rlabel metal2 105644 128681 105644 128681 0 uri_io_oeb\[18\]
rlabel metal2 107660 128709 107660 128709 0 uri_io_oeb\[19\]
rlabel metal2 109676 128765 109676 128765 0 uri_io_oeb\[20\]
rlabel metal2 116844 126567 116844 126567 0 uri_io_oeb\[21\]
rlabel metal2 117516 125895 117516 125895 0 uri_io_oeb\[22\]
rlabel metal2 118188 125811 118188 125811 0 uri_io_oeb\[23\]
rlabel metal3 118300 128884 118300 128884 0 uri_io_oeb\[24\]
rlabel metal2 119637 130060 119637 130060 0 uri_io_oeb\[25\]
rlabel metal2 120204 125951 120204 125951 0 uri_io_oeb\[26\]
rlabel metal2 85484 128233 85484 128233 0 uri_io_oeb\[8\]
rlabel metal2 108780 125727 108780 125727 0 uri_io_oeb\[9\]
rlabel metal2 106820 128744 106820 128744 0 uri_io_out\[10\]
rlabel metal2 92204 128345 92204 128345 0 uri_io_out\[11\]
rlabel metal2 94220 129549 94220 129549 0 uri_io_out\[12\]
rlabel metal2 96236 128373 96236 128373 0 uri_io_out\[13\]
rlabel metal2 98252 129577 98252 129577 0 uri_io_out\[14\]
rlabel metal2 100268 128429 100268 128429 0 uri_io_out\[15\]
rlabel metal2 102284 128653 102284 128653 0 uri_io_out\[16\]
rlabel metal2 104300 128177 104300 128177 0 uri_io_out\[17\]
rlabel metal2 106316 129185 106316 129185 0 uri_io_out\[18\]
rlabel metal2 108332 128737 108332 128737 0 uri_io_out\[19\]
rlabel metal2 116396 125699 116396 125699 0 uri_io_out\[20\]
rlabel metal2 116977 124964 116977 124964 0 uri_io_out\[21\]
rlabel metal2 117740 125783 117740 125783 0 uri_io_out\[22\]
rlabel metal2 118412 125755 118412 125755 0 uri_io_out\[23\]
rlabel metal3 118748 128828 118748 128828 0 uri_io_out\[24\]
rlabel metal2 119756 125923 119756 125923 0 uri_io_out\[25\]
rlabel metal2 120491 124964 120491 124964 0 uri_io_out\[26\]
rlabel metal2 86156 129493 86156 129493 0 uri_io_out\[8\]
rlabel metal2 109004 125755 109004 125755 0 uri_io_out\[9\]
rlabel metal2 83468 128317 83468 128317 0 uri_rst
rlabel metal3 177772 167580 177772 167580 0 vgasp_clk
rlabel metal3 189308 167188 189308 167188 0 vgasp_io_in\[18\]
rlabel metal3 188692 167244 188692 167244 0 vgasp_io_in\[19\]
rlabel metal2 187243 170044 187243 170044 0 vgasp_io_in\[20\]
rlabel metal2 186620 165004 186620 165004 0 vgasp_io_in\[21\]
rlabel metal2 185997 170044 185997 170044 0 vgasp_io_in\[22\]
rlabel metal2 185381 170044 185381 170044 0 vgasp_io_in\[23\]
rlabel metal2 184716 167188 184716 167188 0 vgasp_io_in\[24\]
rlabel metal2 183813 159964 183813 159964 0 vgasp_io_in\[25\]
rlabel metal3 182980 164612 182980 164612 0 vgasp_io_in\[26\]
rlabel metal3 182364 164612 182364 164612 0 vgasp_io_in\[27\]
rlabel metal3 183148 167188 183148 167188 0 vgasp_io_in\[28\]
rlabel metal3 182532 167244 182532 167244 0 vgasp_io_in\[29\]
rlabel metal2 180572 164283 180572 164283 0 vgasp_io_in\[30\]
rlabel metal2 179900 164255 179900 164255 0 vgasp_io_in\[31\]
rlabel metal2 179228 164227 179228 164227 0 vgasp_io_in\[32\]
rlabel metal2 175868 164199 175868 164199 0 vgasp_io_in\[37\]
rlabel metal2 175196 162939 175196 162939 0 vgasp_rst
rlabel metal2 203980 166285 203980 166285 0 vgasp_uio_oe\[0\]
rlabel metal2 203420 166341 203420 166341 0 vgasp_uio_oe\[1\]
rlabel metal2 202860 166369 202860 166369 0 vgasp_uio_oe\[2\]
rlabel metal2 202300 166397 202300 166397 0 vgasp_uio_oe\[3\]
rlabel metal2 201740 166425 201740 166425 0 vgasp_uio_oe\[4\]
rlabel metal2 201180 166453 201180 166453 0 vgasp_uio_oe\[5\]
rlabel metal3 202076 162428 202076 162428 0 vgasp_uio_oe\[6\]
rlabel metal3 201684 162484 201684 162484 0 vgasp_uio_oe\[7\]
rlabel metal2 199500 169393 199500 169393 0 vgasp_uio_out\[0\]
rlabel metal3 200704 162540 200704 162540 0 vgasp_uio_out\[1\]
rlabel metal2 198380 169365 198380 169365 0 vgasp_uio_out\[2\]
rlabel metal2 201180 162372 201180 162372 0 vgasp_uio_out\[3\]
rlabel metal3 202580 168588 202580 168588 0 vgasp_uio_out\[4\]
rlabel metal2 196700 165865 196700 165865 0 vgasp_uio_out\[5\]
rlabel metal3 201796 168420 201796 168420 0 vgasp_uio_out\[6\]
rlabel metal2 195580 165893 195580 165893 0 vgasp_uio_out\[7\]
rlabel metal3 200564 168476 200564 168476 0 vgasp_uo_out\[0\]
rlabel metal2 194460 165921 194460 165921 0 vgasp_uo_out\[1\]
rlabel metal3 199332 168532 199332 168532 0 vgasp_uo_out\[2\]
rlabel metal2 204092 160923 204092 160923 0 vgasp_uo_out\[3\]
rlabel metal2 203420 160951 203420 160951 0 vgasp_uo_out\[4\]
rlabel metal2 192220 166005 192220 166005 0 vgasp_uo_out\[5\]
rlabel metal2 191660 169337 191660 169337 0 vgasp_uo_out\[6\]
rlabel metal2 191100 166033 191100 166033 0 vgasp_uo_out\[7\]
rlabel metal2 5796 1155 5796 1155 0 wb_clk_i
rlabel metal2 6692 1183 6692 1183 0 wb_rst_i
rlabel metal2 7588 3675 7588 3675 0 wbs_ack_o
rlabel metal2 11508 1211 11508 1211 0 wbs_adr_i[0]
rlabel metal2 45500 74081 45500 74081 0 wbs_adr_i[10]
rlabel metal2 46732 1155 46732 1155 0 wbs_adr_i[11]
rlabel metal2 49476 37485 49476 37485 0 wbs_adr_i[12]
rlabel metal3 51940 73108 51940 73108 0 wbs_adr_i[13]
rlabel metal3 54376 73164 54376 73164 0 wbs_adr_i[14]
rlabel metal2 58044 1351 58044 1351 0 wbs_adr_i[15]
rlabel metal3 59248 2100 59248 2100 0 wbs_adr_i[16]
rlabel metal2 59612 38773 59612 38773 0 wbs_adr_i[17]
rlabel metal2 61628 38605 61628 38605 0 wbs_adr_i[18]
rlabel metal2 69468 1155 69468 1155 0 wbs_adr_i[19]
rlabel metal2 15316 1631 15316 1631 0 wbs_adr_i[1]
rlabel metal2 72324 1183 72324 1183 0 wbs_adr_i[20]
rlabel metal2 75180 1239 75180 1239 0 wbs_adr_i[21]
rlabel metal2 69692 39137 69692 39137 0 wbs_adr_i[22]
rlabel metal2 80892 1659 80892 1659 0 wbs_adr_i[23]
rlabel metal2 83748 1603 83748 1603 0 wbs_adr_i[24]
rlabel metal2 86604 1771 86604 1771 0 wbs_adr_i[25]
rlabel metal2 89460 1743 89460 1743 0 wbs_adr_i[26]
rlabel metal3 79996 73108 79996 73108 0 wbs_adr_i[27]
rlabel metal2 95172 1659 95172 1659 0 wbs_adr_i[28]
rlabel metal2 98028 1631 98028 1631 0 wbs_adr_i[29]
rlabel metal2 19124 1155 19124 1155 0 wbs_adr_i[2]
rlabel metal2 85820 39025 85820 39025 0 wbs_adr_i[30]
rlabel metal2 103740 1575 103740 1575 0 wbs_adr_i[31]
rlabel metal2 22932 1183 22932 1183 0 wbs_adr_i[3]
rlabel metal2 26740 1211 26740 1211 0 wbs_adr_i[4]
rlabel metal2 35420 74389 35420 74389 0 wbs_adr_i[5]
rlabel metal2 37436 38689 37436 38689 0 wbs_adr_i[6]
rlabel metal2 35252 1155 35252 1155 0 wbs_adr_i[7]
rlabel metal2 38164 1267 38164 1267 0 wbs_adr_i[8]
rlabel metal2 41020 1183 41020 1183 0 wbs_adr_i[9]
rlabel metal2 8652 1575 8652 1575 0 wbs_cyc_i
rlabel metal2 12460 1603 12460 1603 0 wbs_dat_i[0]
rlabel metal2 46172 38745 46172 38745 0 wbs_dat_i[10]
rlabel metal2 47684 1155 47684 1155 0 wbs_dat_i[11]
rlabel metal2 50316 2100 50316 2100 0 wbs_dat_i[12]
rlabel metal3 52752 73164 52752 73164 0 wbs_dat_i[13]
rlabel metal3 55188 73276 55188 73276 0 wbs_dat_i[14]
rlabel metal2 58996 1211 58996 1211 0 wbs_dat_i[15]
rlabel metal3 60060 2044 60060 2044 0 wbs_dat_i[16]
rlabel metal2 60284 38633 60284 38633 0 wbs_dat_i[17]
rlabel metal2 62300 74333 62300 74333 0 wbs_dat_i[18]
rlabel metal2 70420 1323 70420 1323 0 wbs_dat_i[19]
rlabel metal2 26012 74389 26012 74389 0 wbs_dat_i[1]
rlabel metal2 73276 1267 73276 1267 0 wbs_dat_i[20]
rlabel metal2 72660 37968 72660 37968 0 wbs_dat_i[21]
rlabel metal2 70364 39109 70364 39109 0 wbs_dat_i[22]
rlabel metal2 81844 1631 81844 1631 0 wbs_dat_i[23]
rlabel metal2 74396 74305 74396 74305 0 wbs_dat_i[24]
rlabel metal2 87556 1575 87556 1575 0 wbs_dat_i[25]
rlabel metal2 90412 1211 90412 1211 0 wbs_dat_i[26]
rlabel metal2 93268 1687 93268 1687 0 wbs_dat_i[27]
rlabel metal2 96124 1267 96124 1267 0 wbs_dat_i[28]
rlabel metal2 84476 74473 84476 74473 0 wbs_dat_i[29]
rlabel metal3 22764 2212 22764 2212 0 wbs_dat_i[2]
rlabel metal2 86492 38577 86492 38577 0 wbs_dat_i[30]
rlabel metal3 96740 2324 96740 2324 0 wbs_dat_i[31]
rlabel metal2 23884 1127 23884 1127 0 wbs_dat_i[3]
rlabel metal2 27692 1239 27692 1239 0 wbs_dat_i[4]
rlabel metal2 36092 74277 36092 74277 0 wbs_dat_i[5]
rlabel metal2 38108 38661 38108 38661 0 wbs_dat_i[6]
rlabel metal2 36260 1323 36260 1323 0 wbs_dat_i[7]
rlabel metal2 39004 36855 39004 36855 0 wbs_dat_i[8]
rlabel metal3 43008 73164 43008 73164 0 wbs_dat_i[9]
rlabel metal2 13300 36911 13300 36911 0 wbs_dat_o[0]
rlabel metal2 45780 1183 45780 1183 0 wbs_dat_o[10]
rlabel metal2 48636 73108 48636 73108 0 wbs_dat_o[11]
rlabel metal2 51051 75068 51051 75068 0 wbs_dat_o[12]
rlabel metal3 53536 73108 53536 73108 0 wbs_dat_o[13]
rlabel metal2 57148 36715 57148 36715 0 wbs_dat_o[14]
rlabel metal2 59948 36883 59948 36883 0 wbs_dat_o[15]
rlabel metal3 60872 73108 60872 73108 0 wbs_dat_o[16]
rlabel metal2 60956 38661 60956 38661 0 wbs_dat_o[17]
rlabel metal2 62972 74277 62972 74277 0 wbs_dat_o[18]
rlabel metal3 70364 2044 70364 2044 0 wbs_dat_o[19]
rlabel metal2 26684 39081 26684 39081 0 wbs_dat_o[1]
rlabel metal3 72604 2100 72604 2100 0 wbs_dat_o[20]
rlabel metal3 70896 73108 70896 73108 0 wbs_dat_o[21]
rlabel metal3 72268 73164 72268 73164 0 wbs_dat_o[22]
rlabel metal2 82796 1183 82796 1183 0 wbs_dat_o[23]
rlabel metal2 85708 1155 85708 1155 0 wbs_dat_o[24]
rlabel metal3 88144 2044 88144 2044 0 wbs_dat_o[25]
rlabel metal3 89992 2548 89992 2548 0 wbs_dat_o[26]
rlabel metal3 93940 2156 93940 2156 0 wbs_dat_o[27]
rlabel metal3 97076 2184 97076 2184 0 wbs_dat_o[28]
rlabel metal2 85148 74305 85148 74305 0 wbs_dat_o[29]
rlabel metal2 24892 37744 24892 37744 0 wbs_dat_o[2]
rlabel metal2 97860 37996 97860 37996 0 wbs_dat_o[30]
rlabel metal2 105644 1183 105644 1183 0 wbs_dat_o[31]
rlabel metal2 24836 1211 24836 1211 0 wbs_dat_o[3]
rlabel metal2 34748 74361 34748 74361 0 wbs_dat_o[4]
rlabel metal3 34244 2128 34244 2128 0 wbs_dat_o[5]
rlabel metal2 34356 1155 34356 1155 0 wbs_dat_o[6]
rlabel metal2 37212 1351 37212 1351 0 wbs_dat_o[7]
rlabel metal2 40068 1155 40068 1155 0 wbs_dat_o[8]
rlabel metal2 42924 1155 42924 1155 0 wbs_dat_o[9]
rlabel metal2 14308 36939 14308 36939 0 wbs_sel_i[0]
rlabel metal2 27356 39109 27356 39109 0 wbs_sel_i[1]
rlabel metal2 21868 36855 21868 36855 0 wbs_sel_i[2]
rlabel metal2 25788 1183 25788 1183 0 wbs_sel_i[3]
rlabel metal3 15400 73500 15400 73500 0 wbs_stb_i
rlabel metal2 10444 36883 10444 36883 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 298020 298020
<< end >>
