magic
tech gf180mcuD
magscale 1 5
timestamp 1702301904
<< obsm1 >>
rect 672 463 239288 28545
<< metal2 >>
rect 3360 29600 3416 30000
rect 4032 29600 4088 30000
rect 4704 29600 4760 30000
rect 5376 29600 5432 30000
rect 6048 29600 6104 30000
rect 6720 29600 6776 30000
rect 7392 29600 7448 30000
rect 8064 29600 8120 30000
rect 8736 29600 8792 30000
rect 9408 29600 9464 30000
rect 10080 29600 10136 30000
rect 10752 29600 10808 30000
rect 11424 29600 11480 30000
rect 12096 29600 12152 30000
rect 12768 29600 12824 30000
rect 13440 29600 13496 30000
rect 14112 29600 14168 30000
rect 14784 29600 14840 30000
rect 15456 29600 15512 30000
rect 16128 29600 16184 30000
rect 16800 29600 16856 30000
rect 17472 29600 17528 30000
rect 18144 29600 18200 30000
rect 18816 29600 18872 30000
rect 19488 29600 19544 30000
rect 20160 29600 20216 30000
rect 20832 29600 20888 30000
rect 21504 29600 21560 30000
rect 22176 29600 22232 30000
rect 22848 29600 22904 30000
rect 23520 29600 23576 30000
rect 24192 29600 24248 30000
rect 24864 29600 24920 30000
rect 25536 29600 25592 30000
rect 26208 29600 26264 30000
rect 26880 29600 26936 30000
rect 27552 29600 27608 30000
rect 28224 29600 28280 30000
rect 28896 29600 28952 30000
rect 29568 29600 29624 30000
rect 30240 29600 30296 30000
rect 30912 29600 30968 30000
rect 31584 29600 31640 30000
rect 32256 29600 32312 30000
rect 32928 29600 32984 30000
rect 33600 29600 33656 30000
rect 34272 29600 34328 30000
rect 34944 29600 35000 30000
rect 35616 29600 35672 30000
rect 36288 29600 36344 30000
rect 36960 29600 37016 30000
rect 37632 29600 37688 30000
rect 38304 29600 38360 30000
rect 38976 29600 39032 30000
rect 39648 29600 39704 30000
rect 40320 29600 40376 30000
rect 40992 29600 41048 30000
rect 41664 29600 41720 30000
rect 42336 29600 42392 30000
rect 43008 29600 43064 30000
rect 43680 29600 43736 30000
rect 44352 29600 44408 30000
rect 45024 29600 45080 30000
rect 45696 29600 45752 30000
rect 46368 29600 46424 30000
rect 47040 29600 47096 30000
rect 47712 29600 47768 30000
rect 48384 29600 48440 30000
rect 49056 29600 49112 30000
rect 56448 29600 56504 30000
rect 57120 29600 57176 30000
rect 57792 29600 57848 30000
rect 58464 29600 58520 30000
rect 59136 29600 59192 30000
rect 59808 29600 59864 30000
rect 60480 29600 60536 30000
rect 61152 29600 61208 30000
rect 61824 29600 61880 30000
rect 62496 29600 62552 30000
rect 63168 29600 63224 30000
rect 63840 29600 63896 30000
rect 71232 29600 71288 30000
rect 71904 29600 71960 30000
rect 72576 29600 72632 30000
rect 73248 29600 73304 30000
rect 73920 29600 73976 30000
rect 74592 29600 74648 30000
rect 75264 29600 75320 30000
rect 75936 29600 75992 30000
rect 76608 29600 76664 30000
rect 77280 29600 77336 30000
rect 77952 29600 78008 30000
rect 78624 29600 78680 30000
rect 79296 29600 79352 30000
rect 79968 29600 80024 30000
rect 80640 29600 80696 30000
rect 81312 29600 81368 30000
rect 81984 29600 82040 30000
rect 82656 29600 82712 30000
rect 83328 29600 83384 30000
rect 84000 29600 84056 30000
rect 84672 29600 84728 30000
rect 85344 29600 85400 30000
rect 86016 29600 86072 30000
rect 86688 29600 86744 30000
rect 87360 29600 87416 30000
rect 88032 29600 88088 30000
rect 88704 29600 88760 30000
rect 89376 29600 89432 30000
rect 90048 29600 90104 30000
rect 90720 29600 90776 30000
rect 91392 29600 91448 30000
rect 92064 29600 92120 30000
rect 92736 29600 92792 30000
rect 93408 29600 93464 30000
rect 94080 29600 94136 30000
rect 94752 29600 94808 30000
rect 95424 29600 95480 30000
rect 96096 29600 96152 30000
rect 96768 29600 96824 30000
rect 97440 29600 97496 30000
rect 98112 29600 98168 30000
rect 98784 29600 98840 30000
rect 99456 29600 99512 30000
rect 100128 29600 100184 30000
rect 100800 29600 100856 30000
rect 101472 29600 101528 30000
rect 102144 29600 102200 30000
rect 102816 29600 102872 30000
rect 103488 29600 103544 30000
rect 104160 29600 104216 30000
rect 104832 29600 104888 30000
rect 105504 29600 105560 30000
rect 106176 29600 106232 30000
rect 106848 29600 106904 30000
rect 107520 29600 107576 30000
rect 108192 29600 108248 30000
rect 108864 29600 108920 30000
rect 109536 29600 109592 30000
rect 110208 29600 110264 30000
rect 110880 29600 110936 30000
rect 111552 29600 111608 30000
rect 112224 29600 112280 30000
rect 112896 29600 112952 30000
rect 113568 29600 113624 30000
rect 114240 29600 114296 30000
rect 114912 29600 114968 30000
rect 115584 29600 115640 30000
rect 116256 29600 116312 30000
rect 116928 29600 116984 30000
rect 144480 29600 144536 30000
rect 145152 29600 145208 30000
rect 145824 29600 145880 30000
rect 146496 29600 146552 30000
rect 147168 29600 147224 30000
rect 147840 29600 147896 30000
rect 148512 29600 148568 30000
rect 149184 29600 149240 30000
rect 149856 29600 149912 30000
rect 150528 29600 150584 30000
rect 151200 29600 151256 30000
rect 151872 29600 151928 30000
rect 152544 29600 152600 30000
rect 153216 29600 153272 30000
rect 153888 29600 153944 30000
rect 154560 29600 154616 30000
rect 155232 29600 155288 30000
rect 155904 29600 155960 30000
rect 156576 29600 156632 30000
rect 157248 29600 157304 30000
rect 157920 29600 157976 30000
rect 158592 29600 158648 30000
rect 159264 29600 159320 30000
rect 159936 29600 159992 30000
rect 160608 29600 160664 30000
rect 161280 29600 161336 30000
rect 161952 29600 162008 30000
rect 162624 29600 162680 30000
rect 163296 29600 163352 30000
rect 163968 29600 164024 30000
rect 164640 29600 164696 30000
rect 165312 29600 165368 30000
rect 165984 29600 166040 30000
rect 166656 29600 166712 30000
rect 167328 29600 167384 30000
rect 168000 29600 168056 30000
rect 168672 29600 168728 30000
rect 169344 29600 169400 30000
rect 170016 29600 170072 30000
rect 170688 29600 170744 30000
rect 171360 29600 171416 30000
rect 172032 29600 172088 30000
rect 172704 29600 172760 30000
rect 173376 29600 173432 30000
rect 174048 29600 174104 30000
rect 174720 29600 174776 30000
rect 175392 29600 175448 30000
rect 176064 29600 176120 30000
rect 176736 29600 176792 30000
rect 177408 29600 177464 30000
rect 178080 29600 178136 30000
rect 178752 29600 178808 30000
rect 179424 29600 179480 30000
rect 180096 29600 180152 30000
rect 180768 29600 180824 30000
rect 181440 29600 181496 30000
rect 182112 29600 182168 30000
rect 182784 29600 182840 30000
rect 183456 29600 183512 30000
rect 184128 29600 184184 30000
rect 184800 29600 184856 30000
rect 185472 29600 185528 30000
rect 186144 29600 186200 30000
rect 186816 29600 186872 30000
rect 190848 29600 190904 30000
rect 191520 29600 191576 30000
rect 192192 29600 192248 30000
rect 192864 29600 192920 30000
rect 193536 29600 193592 30000
rect 194208 29600 194264 30000
rect 194880 29600 194936 30000
rect 195552 29600 195608 30000
rect 196224 29600 196280 30000
rect 200256 29600 200312 30000
rect 200928 29600 200984 30000
rect 201600 29600 201656 30000
rect 202272 29600 202328 30000
rect 202944 29600 203000 30000
rect 203616 29600 203672 30000
rect 204288 29600 204344 30000
rect 204960 29600 205016 30000
rect 205632 29600 205688 30000
rect 206304 29600 206360 30000
rect 206976 29600 207032 30000
rect 207648 29600 207704 30000
rect 208320 29600 208376 30000
rect 208992 29600 209048 30000
rect 209664 29600 209720 30000
rect 210336 29600 210392 30000
rect 211008 29600 211064 30000
rect 211680 29600 211736 30000
rect 212352 29600 212408 30000
rect 213024 29600 213080 30000
rect 213696 29600 213752 30000
rect 214368 29600 214424 30000
rect 215040 29600 215096 30000
rect 215712 29600 215768 30000
rect 216384 29600 216440 30000
rect 217056 29600 217112 30000
rect 217728 29600 217784 30000
rect 218400 29600 218456 30000
rect 219072 29600 219128 30000
rect 219744 29600 219800 30000
rect 220416 29600 220472 30000
rect 221088 29600 221144 30000
rect 221760 29600 221816 30000
rect 222432 29600 222488 30000
rect 223104 29600 223160 30000
rect 223776 29600 223832 30000
rect 224448 29600 224504 30000
rect 225120 29600 225176 30000
rect 225792 29600 225848 30000
rect 226464 29600 226520 30000
rect 227136 29600 227192 30000
rect 227808 29600 227864 30000
rect 228480 29600 228536 30000
rect 229152 29600 229208 30000
rect 229824 29600 229880 30000
rect 230496 29600 230552 30000
rect 231168 29600 231224 30000
rect 231840 29600 231896 30000
rect 232512 29600 232568 30000
rect 233184 29600 233240 30000
rect 233856 29600 233912 30000
rect 234528 29600 234584 30000
rect 235200 29600 235256 30000
rect 235872 29600 235928 30000
rect 236544 29600 236600 30000
rect 4368 0 4424 400
rect 5040 0 5096 400
rect 5712 0 5768 400
rect 6384 0 6440 400
rect 7056 0 7112 400
rect 7728 0 7784 400
rect 8400 0 8456 400
rect 9072 0 9128 400
rect 9744 0 9800 400
rect 10416 0 10472 400
rect 11088 0 11144 400
rect 11760 0 11816 400
rect 12432 0 12488 400
rect 13104 0 13160 400
rect 13776 0 13832 400
rect 14448 0 14504 400
rect 15120 0 15176 400
rect 15792 0 15848 400
rect 16464 0 16520 400
rect 17136 0 17192 400
rect 17808 0 17864 400
rect 18480 0 18536 400
rect 19152 0 19208 400
rect 19824 0 19880 400
rect 20496 0 20552 400
rect 21168 0 21224 400
rect 21840 0 21896 400
rect 22512 0 22568 400
rect 23184 0 23240 400
rect 23856 0 23912 400
rect 24528 0 24584 400
rect 25200 0 25256 400
rect 25872 0 25928 400
rect 26544 0 26600 400
rect 27216 0 27272 400
rect 27888 0 27944 400
rect 28560 0 28616 400
rect 29232 0 29288 400
rect 29904 0 29960 400
rect 30576 0 30632 400
rect 31248 0 31304 400
rect 31920 0 31976 400
rect 32592 0 32648 400
rect 33264 0 33320 400
rect 33936 0 33992 400
rect 34608 0 34664 400
rect 35280 0 35336 400
rect 35952 0 36008 400
rect 36624 0 36680 400
rect 37296 0 37352 400
rect 37968 0 38024 400
rect 38640 0 38696 400
rect 39312 0 39368 400
rect 39984 0 40040 400
rect 40656 0 40712 400
rect 41328 0 41384 400
rect 42000 0 42056 400
rect 42672 0 42728 400
rect 43344 0 43400 400
rect 44016 0 44072 400
rect 44688 0 44744 400
rect 45360 0 45416 400
rect 46032 0 46088 400
rect 46704 0 46760 400
rect 47376 0 47432 400
rect 48048 0 48104 400
rect 48720 0 48776 400
rect 52752 0 52808 400
rect 53424 0 53480 400
rect 54096 0 54152 400
rect 54768 0 54824 400
rect 55440 0 55496 400
rect 56112 0 56168 400
rect 56784 0 56840 400
rect 57456 0 57512 400
rect 58128 0 58184 400
rect 58800 0 58856 400
rect 59472 0 59528 400
rect 60144 0 60200 400
rect 60816 0 60872 400
rect 61488 0 61544 400
rect 62160 0 62216 400
rect 62832 0 62888 400
rect 63504 0 63560 400
rect 64176 0 64232 400
rect 64848 0 64904 400
rect 65520 0 65576 400
rect 66192 0 66248 400
rect 66864 0 66920 400
rect 67536 0 67592 400
rect 68208 0 68264 400
rect 68880 0 68936 400
rect 69552 0 69608 400
rect 70224 0 70280 400
rect 70896 0 70952 400
rect 71568 0 71624 400
rect 72240 0 72296 400
rect 72912 0 72968 400
rect 73584 0 73640 400
rect 74256 0 74312 400
rect 74928 0 74984 400
rect 75600 0 75656 400
rect 76272 0 76328 400
rect 76944 0 77000 400
rect 77616 0 77672 400
rect 78288 0 78344 400
rect 78960 0 79016 400
rect 79632 0 79688 400
rect 80304 0 80360 400
rect 80976 0 81032 400
rect 81648 0 81704 400
rect 82320 0 82376 400
rect 82992 0 83048 400
rect 83664 0 83720 400
rect 84336 0 84392 400
rect 85008 0 85064 400
rect 85680 0 85736 400
rect 86352 0 86408 400
rect 87024 0 87080 400
rect 87696 0 87752 400
rect 88368 0 88424 400
rect 89040 0 89096 400
rect 89712 0 89768 400
rect 90384 0 90440 400
rect 91056 0 91112 400
rect 91728 0 91784 400
rect 92400 0 92456 400
rect 93072 0 93128 400
rect 93744 0 93800 400
rect 94416 0 94472 400
rect 95088 0 95144 400
rect 95760 0 95816 400
rect 96432 0 96488 400
rect 97104 0 97160 400
rect 97776 0 97832 400
rect 98448 0 98504 400
rect 99120 0 99176 400
rect 99792 0 99848 400
rect 100464 0 100520 400
rect 101136 0 101192 400
rect 101808 0 101864 400
rect 102480 0 102536 400
rect 103152 0 103208 400
rect 103824 0 103880 400
rect 104496 0 104552 400
rect 105168 0 105224 400
rect 112560 0 112616 400
rect 113232 0 113288 400
rect 113904 0 113960 400
rect 114576 0 114632 400
rect 115248 0 115304 400
rect 115920 0 115976 400
rect 116592 0 116648 400
rect 117264 0 117320 400
rect 117936 0 117992 400
rect 118608 0 118664 400
rect 119280 0 119336 400
rect 119952 0 120008 400
rect 120624 0 120680 400
rect 121296 0 121352 400
rect 121968 0 122024 400
rect 122640 0 122696 400
rect 143472 0 143528 400
rect 144144 0 144200 400
rect 144816 0 144872 400
rect 145488 0 145544 400
rect 146160 0 146216 400
rect 146832 0 146888 400
rect 147504 0 147560 400
rect 148176 0 148232 400
rect 148848 0 148904 400
rect 149520 0 149576 400
rect 150192 0 150248 400
rect 150864 0 150920 400
rect 151536 0 151592 400
rect 152208 0 152264 400
rect 152880 0 152936 400
rect 153552 0 153608 400
rect 154224 0 154280 400
rect 154896 0 154952 400
rect 155568 0 155624 400
rect 156240 0 156296 400
rect 156912 0 156968 400
rect 157584 0 157640 400
rect 158256 0 158312 400
rect 158928 0 158984 400
rect 159600 0 159656 400
rect 160272 0 160328 400
rect 160944 0 161000 400
rect 161616 0 161672 400
rect 162288 0 162344 400
rect 162960 0 163016 400
rect 163632 0 163688 400
rect 164304 0 164360 400
rect 164976 0 165032 400
rect 165648 0 165704 400
rect 166320 0 166376 400
rect 166992 0 167048 400
rect 167664 0 167720 400
rect 168336 0 168392 400
rect 169008 0 169064 400
rect 169680 0 169736 400
rect 170352 0 170408 400
rect 171024 0 171080 400
rect 171696 0 171752 400
rect 172368 0 172424 400
rect 173040 0 173096 400
rect 173712 0 173768 400
rect 174384 0 174440 400
rect 175056 0 175112 400
rect 175728 0 175784 400
rect 176400 0 176456 400
rect 177072 0 177128 400
rect 177744 0 177800 400
rect 178416 0 178472 400
rect 179088 0 179144 400
rect 179760 0 179816 400
rect 180432 0 180488 400
rect 181104 0 181160 400
rect 181776 0 181832 400
rect 182448 0 182504 400
rect 183120 0 183176 400
rect 183792 0 183848 400
rect 184464 0 184520 400
rect 185136 0 185192 400
rect 185808 0 185864 400
rect 186480 0 186536 400
rect 187152 0 187208 400
rect 187824 0 187880 400
rect 188496 0 188552 400
rect 189168 0 189224 400
rect 189840 0 189896 400
rect 190512 0 190568 400
rect 191184 0 191240 400
rect 191856 0 191912 400
rect 192528 0 192584 400
rect 193200 0 193256 400
rect 193872 0 193928 400
rect 194544 0 194600 400
rect 195216 0 195272 400
rect 195888 0 195944 400
rect 196560 0 196616 400
rect 197232 0 197288 400
rect 197904 0 197960 400
rect 198576 0 198632 400
rect 199248 0 199304 400
rect 199920 0 199976 400
rect 200592 0 200648 400
rect 201264 0 201320 400
rect 201936 0 201992 400
rect 202608 0 202664 400
rect 203280 0 203336 400
rect 203952 0 204008 400
rect 204624 0 204680 400
rect 205296 0 205352 400
rect 205968 0 206024 400
rect 206640 0 206696 400
rect 207312 0 207368 400
rect 207984 0 208040 400
rect 208656 0 208712 400
rect 209328 0 209384 400
rect 210000 0 210056 400
rect 210672 0 210728 400
rect 211344 0 211400 400
rect 212016 0 212072 400
rect 212688 0 212744 400
rect 213360 0 213416 400
<< obsm2 >>
rect 854 29570 3330 29666
rect 3446 29570 4002 29666
rect 4118 29570 4674 29666
rect 4790 29570 5346 29666
rect 5462 29570 6018 29666
rect 6134 29570 6690 29666
rect 6806 29570 7362 29666
rect 7478 29570 8034 29666
rect 8150 29570 8706 29666
rect 8822 29570 9378 29666
rect 9494 29570 10050 29666
rect 10166 29570 10722 29666
rect 10838 29570 11394 29666
rect 11510 29570 12066 29666
rect 12182 29570 12738 29666
rect 12854 29570 13410 29666
rect 13526 29570 14082 29666
rect 14198 29570 14754 29666
rect 14870 29570 15426 29666
rect 15542 29570 16098 29666
rect 16214 29570 16770 29666
rect 16886 29570 17442 29666
rect 17558 29570 18114 29666
rect 18230 29570 18786 29666
rect 18902 29570 19458 29666
rect 19574 29570 20130 29666
rect 20246 29570 20802 29666
rect 20918 29570 21474 29666
rect 21590 29570 22146 29666
rect 22262 29570 22818 29666
rect 22934 29570 23490 29666
rect 23606 29570 24162 29666
rect 24278 29570 24834 29666
rect 24950 29570 25506 29666
rect 25622 29570 26178 29666
rect 26294 29570 26850 29666
rect 26966 29570 27522 29666
rect 27638 29570 28194 29666
rect 28310 29570 28866 29666
rect 28982 29570 29538 29666
rect 29654 29570 30210 29666
rect 30326 29570 30882 29666
rect 30998 29570 31554 29666
rect 31670 29570 32226 29666
rect 32342 29570 32898 29666
rect 33014 29570 33570 29666
rect 33686 29570 34242 29666
rect 34358 29570 34914 29666
rect 35030 29570 35586 29666
rect 35702 29570 36258 29666
rect 36374 29570 36930 29666
rect 37046 29570 37602 29666
rect 37718 29570 38274 29666
rect 38390 29570 38946 29666
rect 39062 29570 39618 29666
rect 39734 29570 40290 29666
rect 40406 29570 40962 29666
rect 41078 29570 41634 29666
rect 41750 29570 42306 29666
rect 42422 29570 42978 29666
rect 43094 29570 43650 29666
rect 43766 29570 44322 29666
rect 44438 29570 44994 29666
rect 45110 29570 45666 29666
rect 45782 29570 46338 29666
rect 46454 29570 47010 29666
rect 47126 29570 47682 29666
rect 47798 29570 48354 29666
rect 48470 29570 49026 29666
rect 49142 29570 56418 29666
rect 56534 29570 57090 29666
rect 57206 29570 57762 29666
rect 57878 29570 58434 29666
rect 58550 29570 59106 29666
rect 59222 29570 59778 29666
rect 59894 29570 60450 29666
rect 60566 29570 61122 29666
rect 61238 29570 61794 29666
rect 61910 29570 62466 29666
rect 62582 29570 63138 29666
rect 63254 29570 63810 29666
rect 63926 29570 71202 29666
rect 71318 29570 71874 29666
rect 71990 29570 72546 29666
rect 72662 29570 73218 29666
rect 73334 29570 73890 29666
rect 74006 29570 74562 29666
rect 74678 29570 75234 29666
rect 75350 29570 75906 29666
rect 76022 29570 76578 29666
rect 76694 29570 77250 29666
rect 77366 29570 77922 29666
rect 78038 29570 78594 29666
rect 78710 29570 79266 29666
rect 79382 29570 79938 29666
rect 80054 29570 80610 29666
rect 80726 29570 81282 29666
rect 81398 29570 81954 29666
rect 82070 29570 82626 29666
rect 82742 29570 83298 29666
rect 83414 29570 83970 29666
rect 84086 29570 84642 29666
rect 84758 29570 85314 29666
rect 85430 29570 85986 29666
rect 86102 29570 86658 29666
rect 86774 29570 87330 29666
rect 87446 29570 88002 29666
rect 88118 29570 88674 29666
rect 88790 29570 89346 29666
rect 89462 29570 90018 29666
rect 90134 29570 90690 29666
rect 90806 29570 91362 29666
rect 91478 29570 92034 29666
rect 92150 29570 92706 29666
rect 92822 29570 93378 29666
rect 93494 29570 94050 29666
rect 94166 29570 94722 29666
rect 94838 29570 95394 29666
rect 95510 29570 96066 29666
rect 96182 29570 96738 29666
rect 96854 29570 97410 29666
rect 97526 29570 98082 29666
rect 98198 29570 98754 29666
rect 98870 29570 99426 29666
rect 99542 29570 100098 29666
rect 100214 29570 100770 29666
rect 100886 29570 101442 29666
rect 101558 29570 102114 29666
rect 102230 29570 102786 29666
rect 102902 29570 103458 29666
rect 103574 29570 104130 29666
rect 104246 29570 104802 29666
rect 104918 29570 105474 29666
rect 105590 29570 106146 29666
rect 106262 29570 106818 29666
rect 106934 29570 107490 29666
rect 107606 29570 108162 29666
rect 108278 29570 108834 29666
rect 108950 29570 109506 29666
rect 109622 29570 110178 29666
rect 110294 29570 110850 29666
rect 110966 29570 111522 29666
rect 111638 29570 112194 29666
rect 112310 29570 112866 29666
rect 112982 29570 113538 29666
rect 113654 29570 114210 29666
rect 114326 29570 114882 29666
rect 114998 29570 115554 29666
rect 115670 29570 116226 29666
rect 116342 29570 116898 29666
rect 117014 29570 144450 29666
rect 144566 29570 145122 29666
rect 145238 29570 145794 29666
rect 145910 29570 146466 29666
rect 146582 29570 147138 29666
rect 147254 29570 147810 29666
rect 147926 29570 148482 29666
rect 148598 29570 149154 29666
rect 149270 29570 149826 29666
rect 149942 29570 150498 29666
rect 150614 29570 151170 29666
rect 151286 29570 151842 29666
rect 151958 29570 152514 29666
rect 152630 29570 153186 29666
rect 153302 29570 153858 29666
rect 153974 29570 154530 29666
rect 154646 29570 155202 29666
rect 155318 29570 155874 29666
rect 155990 29570 156546 29666
rect 156662 29570 157218 29666
rect 157334 29570 157890 29666
rect 158006 29570 158562 29666
rect 158678 29570 159234 29666
rect 159350 29570 159906 29666
rect 160022 29570 160578 29666
rect 160694 29570 161250 29666
rect 161366 29570 161922 29666
rect 162038 29570 162594 29666
rect 162710 29570 163266 29666
rect 163382 29570 163938 29666
rect 164054 29570 164610 29666
rect 164726 29570 165282 29666
rect 165398 29570 165954 29666
rect 166070 29570 166626 29666
rect 166742 29570 167298 29666
rect 167414 29570 167970 29666
rect 168086 29570 168642 29666
rect 168758 29570 169314 29666
rect 169430 29570 169986 29666
rect 170102 29570 170658 29666
rect 170774 29570 171330 29666
rect 171446 29570 172002 29666
rect 172118 29570 172674 29666
rect 172790 29570 173346 29666
rect 173462 29570 174018 29666
rect 174134 29570 174690 29666
rect 174806 29570 175362 29666
rect 175478 29570 176034 29666
rect 176150 29570 176706 29666
rect 176822 29570 177378 29666
rect 177494 29570 178050 29666
rect 178166 29570 178722 29666
rect 178838 29570 179394 29666
rect 179510 29570 180066 29666
rect 180182 29570 180738 29666
rect 180854 29570 181410 29666
rect 181526 29570 182082 29666
rect 182198 29570 182754 29666
rect 182870 29570 183426 29666
rect 183542 29570 184098 29666
rect 184214 29570 184770 29666
rect 184886 29570 185442 29666
rect 185558 29570 186114 29666
rect 186230 29570 186786 29666
rect 186902 29570 190818 29666
rect 190934 29570 191490 29666
rect 191606 29570 192162 29666
rect 192278 29570 192834 29666
rect 192950 29570 193506 29666
rect 193622 29570 194178 29666
rect 194294 29570 194850 29666
rect 194966 29570 195522 29666
rect 195638 29570 196194 29666
rect 196310 29570 200226 29666
rect 200342 29570 200898 29666
rect 201014 29570 201570 29666
rect 201686 29570 202242 29666
rect 202358 29570 202914 29666
rect 203030 29570 203586 29666
rect 203702 29570 204258 29666
rect 204374 29570 204930 29666
rect 205046 29570 205602 29666
rect 205718 29570 206274 29666
rect 206390 29570 206946 29666
rect 207062 29570 207618 29666
rect 207734 29570 208290 29666
rect 208406 29570 208962 29666
rect 209078 29570 209634 29666
rect 209750 29570 210306 29666
rect 210422 29570 210978 29666
rect 211094 29570 211650 29666
rect 211766 29570 212322 29666
rect 212438 29570 212994 29666
rect 213110 29570 213666 29666
rect 213782 29570 214338 29666
rect 214454 29570 215010 29666
rect 215126 29570 215682 29666
rect 215798 29570 216354 29666
rect 216470 29570 217026 29666
rect 217142 29570 217698 29666
rect 217814 29570 218370 29666
rect 218486 29570 219042 29666
rect 219158 29570 219714 29666
rect 219830 29570 220386 29666
rect 220502 29570 221058 29666
rect 221174 29570 221730 29666
rect 221846 29570 222402 29666
rect 222518 29570 223074 29666
rect 223190 29570 223746 29666
rect 223862 29570 224418 29666
rect 224534 29570 225090 29666
rect 225206 29570 225762 29666
rect 225878 29570 226434 29666
rect 226550 29570 227106 29666
rect 227222 29570 227778 29666
rect 227894 29570 228450 29666
rect 228566 29570 229122 29666
rect 229238 29570 229794 29666
rect 229910 29570 230466 29666
rect 230582 29570 231138 29666
rect 231254 29570 231810 29666
rect 231926 29570 232482 29666
rect 232598 29570 233154 29666
rect 233270 29570 233826 29666
rect 233942 29570 234498 29666
rect 234614 29570 235170 29666
rect 235286 29570 235842 29666
rect 235958 29570 236514 29666
rect 236630 29570 239162 29666
rect 854 430 239162 29570
rect 854 233 4338 430
rect 4454 233 5010 430
rect 5126 233 5682 430
rect 5798 233 6354 430
rect 6470 233 7026 430
rect 7142 233 7698 430
rect 7814 233 8370 430
rect 8486 233 9042 430
rect 9158 233 9714 430
rect 9830 233 10386 430
rect 10502 233 11058 430
rect 11174 233 11730 430
rect 11846 233 12402 430
rect 12518 233 13074 430
rect 13190 233 13746 430
rect 13862 233 14418 430
rect 14534 233 15090 430
rect 15206 233 15762 430
rect 15878 233 16434 430
rect 16550 233 17106 430
rect 17222 233 17778 430
rect 17894 233 18450 430
rect 18566 233 19122 430
rect 19238 233 19794 430
rect 19910 233 20466 430
rect 20582 233 21138 430
rect 21254 233 21810 430
rect 21926 233 22482 430
rect 22598 233 23154 430
rect 23270 233 23826 430
rect 23942 233 24498 430
rect 24614 233 25170 430
rect 25286 233 25842 430
rect 25958 233 26514 430
rect 26630 233 27186 430
rect 27302 233 27858 430
rect 27974 233 28530 430
rect 28646 233 29202 430
rect 29318 233 29874 430
rect 29990 233 30546 430
rect 30662 233 31218 430
rect 31334 233 31890 430
rect 32006 233 32562 430
rect 32678 233 33234 430
rect 33350 233 33906 430
rect 34022 233 34578 430
rect 34694 233 35250 430
rect 35366 233 35922 430
rect 36038 233 36594 430
rect 36710 233 37266 430
rect 37382 233 37938 430
rect 38054 233 38610 430
rect 38726 233 39282 430
rect 39398 233 39954 430
rect 40070 233 40626 430
rect 40742 233 41298 430
rect 41414 233 41970 430
rect 42086 233 42642 430
rect 42758 233 43314 430
rect 43430 233 43986 430
rect 44102 233 44658 430
rect 44774 233 45330 430
rect 45446 233 46002 430
rect 46118 233 46674 430
rect 46790 233 47346 430
rect 47462 233 48018 430
rect 48134 233 48690 430
rect 48806 233 52722 430
rect 52838 233 53394 430
rect 53510 233 54066 430
rect 54182 233 54738 430
rect 54854 233 55410 430
rect 55526 233 56082 430
rect 56198 233 56754 430
rect 56870 233 57426 430
rect 57542 233 58098 430
rect 58214 233 58770 430
rect 58886 233 59442 430
rect 59558 233 60114 430
rect 60230 233 60786 430
rect 60902 233 61458 430
rect 61574 233 62130 430
rect 62246 233 62802 430
rect 62918 233 63474 430
rect 63590 233 64146 430
rect 64262 233 64818 430
rect 64934 233 65490 430
rect 65606 233 66162 430
rect 66278 233 66834 430
rect 66950 233 67506 430
rect 67622 233 68178 430
rect 68294 233 68850 430
rect 68966 233 69522 430
rect 69638 233 70194 430
rect 70310 233 70866 430
rect 70982 233 71538 430
rect 71654 233 72210 430
rect 72326 233 72882 430
rect 72998 233 73554 430
rect 73670 233 74226 430
rect 74342 233 74898 430
rect 75014 233 75570 430
rect 75686 233 76242 430
rect 76358 233 76914 430
rect 77030 233 77586 430
rect 77702 233 78258 430
rect 78374 233 78930 430
rect 79046 233 79602 430
rect 79718 233 80274 430
rect 80390 233 80946 430
rect 81062 233 81618 430
rect 81734 233 82290 430
rect 82406 233 82962 430
rect 83078 233 83634 430
rect 83750 233 84306 430
rect 84422 233 84978 430
rect 85094 233 85650 430
rect 85766 233 86322 430
rect 86438 233 86994 430
rect 87110 233 87666 430
rect 87782 233 88338 430
rect 88454 233 89010 430
rect 89126 233 89682 430
rect 89798 233 90354 430
rect 90470 233 91026 430
rect 91142 233 91698 430
rect 91814 233 92370 430
rect 92486 233 93042 430
rect 93158 233 93714 430
rect 93830 233 94386 430
rect 94502 233 95058 430
rect 95174 233 95730 430
rect 95846 233 96402 430
rect 96518 233 97074 430
rect 97190 233 97746 430
rect 97862 233 98418 430
rect 98534 233 99090 430
rect 99206 233 99762 430
rect 99878 233 100434 430
rect 100550 233 101106 430
rect 101222 233 101778 430
rect 101894 233 102450 430
rect 102566 233 103122 430
rect 103238 233 103794 430
rect 103910 233 104466 430
rect 104582 233 105138 430
rect 105254 233 112530 430
rect 112646 233 113202 430
rect 113318 233 113874 430
rect 113990 233 114546 430
rect 114662 233 115218 430
rect 115334 233 115890 430
rect 116006 233 116562 430
rect 116678 233 117234 430
rect 117350 233 117906 430
rect 118022 233 118578 430
rect 118694 233 119250 430
rect 119366 233 119922 430
rect 120038 233 120594 430
rect 120710 233 121266 430
rect 121382 233 121938 430
rect 122054 233 122610 430
rect 122726 233 143442 430
rect 143558 233 144114 430
rect 144230 233 144786 430
rect 144902 233 145458 430
rect 145574 233 146130 430
rect 146246 233 146802 430
rect 146918 233 147474 430
rect 147590 233 148146 430
rect 148262 233 148818 430
rect 148934 233 149490 430
rect 149606 233 150162 430
rect 150278 233 150834 430
rect 150950 233 151506 430
rect 151622 233 152178 430
rect 152294 233 152850 430
rect 152966 233 153522 430
rect 153638 233 154194 430
rect 154310 233 154866 430
rect 154982 233 155538 430
rect 155654 233 156210 430
rect 156326 233 156882 430
rect 156998 233 157554 430
rect 157670 233 158226 430
rect 158342 233 158898 430
rect 159014 233 159570 430
rect 159686 233 160242 430
rect 160358 233 160914 430
rect 161030 233 161586 430
rect 161702 233 162258 430
rect 162374 233 162930 430
rect 163046 233 163602 430
rect 163718 233 164274 430
rect 164390 233 164946 430
rect 165062 233 165618 430
rect 165734 233 166290 430
rect 166406 233 166962 430
rect 167078 233 167634 430
rect 167750 233 168306 430
rect 168422 233 168978 430
rect 169094 233 169650 430
rect 169766 233 170322 430
rect 170438 233 170994 430
rect 171110 233 171666 430
rect 171782 233 172338 430
rect 172454 233 173010 430
rect 173126 233 173682 430
rect 173798 233 174354 430
rect 174470 233 175026 430
rect 175142 233 175698 430
rect 175814 233 176370 430
rect 176486 233 177042 430
rect 177158 233 177714 430
rect 177830 233 178386 430
rect 178502 233 179058 430
rect 179174 233 179730 430
rect 179846 233 180402 430
rect 180518 233 181074 430
rect 181190 233 181746 430
rect 181862 233 182418 430
rect 182534 233 183090 430
rect 183206 233 183762 430
rect 183878 233 184434 430
rect 184550 233 185106 430
rect 185222 233 185778 430
rect 185894 233 186450 430
rect 186566 233 187122 430
rect 187238 233 187794 430
rect 187910 233 188466 430
rect 188582 233 189138 430
rect 189254 233 189810 430
rect 189926 233 190482 430
rect 190598 233 191154 430
rect 191270 233 191826 430
rect 191942 233 192498 430
rect 192614 233 193170 430
rect 193286 233 193842 430
rect 193958 233 194514 430
rect 194630 233 195186 430
rect 195302 233 195858 430
rect 195974 233 196530 430
rect 196646 233 197202 430
rect 197318 233 197874 430
rect 197990 233 198546 430
rect 198662 233 199218 430
rect 199334 233 199890 430
rect 200006 233 200562 430
rect 200678 233 201234 430
rect 201350 233 201906 430
rect 202022 233 202578 430
rect 202694 233 203250 430
rect 203366 233 203922 430
rect 204038 233 204594 430
rect 204710 233 205266 430
rect 205382 233 205938 430
rect 206054 233 206610 430
rect 206726 233 207282 430
rect 207398 233 207954 430
rect 208070 233 208626 430
rect 208742 233 209298 430
rect 209414 233 209970 430
rect 210086 233 210642 430
rect 210758 233 211314 430
rect 211430 233 211986 430
rect 212102 233 212658 430
rect 212774 233 213330 430
rect 213446 233 239162 430
<< metal3 >>
rect 239600 29008 240000 29064
rect 239600 28560 240000 28616
rect 239600 28112 240000 28168
rect 0 27776 400 27832
rect 239600 27664 240000 27720
rect 0 27216 400 27272
rect 239600 27216 240000 27272
rect 239600 26768 240000 26824
rect 0 26656 400 26712
rect 239600 26320 240000 26376
rect 0 26096 400 26152
rect 239600 25872 240000 25928
rect 0 25536 400 25592
rect 239600 25424 240000 25480
rect 0 24976 400 25032
rect 239600 24976 240000 25032
rect 239600 24528 240000 24584
rect 0 24416 400 24472
rect 239600 24080 240000 24136
rect 0 23856 400 23912
rect 239600 23632 240000 23688
rect 0 23296 400 23352
rect 239600 23184 240000 23240
rect 0 22736 400 22792
rect 239600 22736 240000 22792
rect 239600 22288 240000 22344
rect 0 22176 400 22232
rect 239600 21840 240000 21896
rect 0 21616 400 21672
rect 239600 21392 240000 21448
rect 0 21056 400 21112
rect 239600 20944 240000 21000
rect 0 20496 400 20552
rect 239600 20496 240000 20552
rect 239600 20048 240000 20104
rect 0 19936 400 19992
rect 239600 19600 240000 19656
rect 0 19376 400 19432
rect 239600 19152 240000 19208
rect 0 18816 400 18872
rect 239600 18704 240000 18760
rect 0 18256 400 18312
rect 239600 18256 240000 18312
rect 239600 17808 240000 17864
rect 0 17696 400 17752
rect 239600 17360 240000 17416
rect 0 17136 400 17192
rect 239600 16912 240000 16968
rect 0 16576 400 16632
rect 239600 16464 240000 16520
rect 0 16016 400 16072
rect 239600 16016 240000 16072
rect 239600 15568 240000 15624
rect 0 15456 400 15512
rect 239600 15120 240000 15176
rect 0 14896 400 14952
rect 239600 14672 240000 14728
rect 0 14336 400 14392
rect 239600 14224 240000 14280
rect 0 13776 400 13832
rect 239600 13776 240000 13832
rect 239600 13328 240000 13384
rect 0 13216 400 13272
rect 239600 12880 240000 12936
rect 0 12656 400 12712
rect 239600 12432 240000 12488
rect 0 12096 400 12152
rect 239600 11984 240000 12040
rect 0 11536 400 11592
rect 239600 11536 240000 11592
rect 239600 11088 240000 11144
rect 0 10976 400 11032
rect 239600 10640 240000 10696
rect 0 10416 400 10472
rect 239600 10192 240000 10248
rect 0 9856 400 9912
rect 239600 9744 240000 9800
rect 0 9296 400 9352
rect 239600 9296 240000 9352
rect 239600 8848 240000 8904
rect 0 8736 400 8792
rect 239600 8400 240000 8456
rect 0 8176 400 8232
rect 239600 7952 240000 8008
rect 0 7616 400 7672
rect 239600 7504 240000 7560
rect 0 7056 400 7112
rect 239600 7056 240000 7112
rect 239600 6608 240000 6664
rect 0 6496 400 6552
rect 239600 6160 240000 6216
rect 0 5936 400 5992
rect 239600 5712 240000 5768
rect 0 5376 400 5432
rect 239600 5264 240000 5320
rect 0 4816 400 4872
rect 239600 4816 240000 4872
rect 239600 4368 240000 4424
rect 0 4256 400 4312
rect 239600 3920 240000 3976
rect 0 3696 400 3752
rect 239600 3472 240000 3528
rect 0 3136 400 3192
rect 239600 3024 240000 3080
rect 0 2576 400 2632
rect 239600 2576 240000 2632
rect 239600 2128 240000 2184
rect 0 2016 400 2072
rect 239600 1680 240000 1736
rect 239600 1232 240000 1288
rect 239600 784 240000 840
<< obsm3 >>
rect 400 28978 239570 29050
rect 400 28646 239666 28978
rect 400 28530 239570 28646
rect 400 28198 239666 28530
rect 400 28082 239570 28198
rect 400 27862 239666 28082
rect 430 27750 239666 27862
rect 430 27746 239570 27750
rect 400 27634 239570 27746
rect 400 27302 239666 27634
rect 430 27186 239570 27302
rect 400 26854 239666 27186
rect 400 26742 239570 26854
rect 430 26738 239570 26742
rect 430 26626 239666 26738
rect 400 26406 239666 26626
rect 400 26290 239570 26406
rect 400 26182 239666 26290
rect 430 26066 239666 26182
rect 400 25958 239666 26066
rect 400 25842 239570 25958
rect 400 25622 239666 25842
rect 430 25510 239666 25622
rect 430 25506 239570 25510
rect 400 25394 239570 25506
rect 400 25062 239666 25394
rect 430 24946 239570 25062
rect 400 24614 239666 24946
rect 400 24502 239570 24614
rect 430 24498 239570 24502
rect 430 24386 239666 24498
rect 400 24166 239666 24386
rect 400 24050 239570 24166
rect 400 23942 239666 24050
rect 430 23826 239666 23942
rect 400 23718 239666 23826
rect 400 23602 239570 23718
rect 400 23382 239666 23602
rect 430 23270 239666 23382
rect 430 23266 239570 23270
rect 400 23154 239570 23266
rect 400 22822 239666 23154
rect 430 22706 239570 22822
rect 400 22374 239666 22706
rect 400 22262 239570 22374
rect 430 22258 239570 22262
rect 430 22146 239666 22258
rect 400 21926 239666 22146
rect 400 21810 239570 21926
rect 400 21702 239666 21810
rect 430 21586 239666 21702
rect 400 21478 239666 21586
rect 400 21362 239570 21478
rect 400 21142 239666 21362
rect 430 21030 239666 21142
rect 430 21026 239570 21030
rect 400 20914 239570 21026
rect 400 20582 239666 20914
rect 430 20466 239570 20582
rect 400 20134 239666 20466
rect 400 20022 239570 20134
rect 430 20018 239570 20022
rect 430 19906 239666 20018
rect 400 19686 239666 19906
rect 400 19570 239570 19686
rect 400 19462 239666 19570
rect 430 19346 239666 19462
rect 400 19238 239666 19346
rect 400 19122 239570 19238
rect 400 18902 239666 19122
rect 430 18790 239666 18902
rect 430 18786 239570 18790
rect 400 18674 239570 18786
rect 400 18342 239666 18674
rect 430 18226 239570 18342
rect 400 17894 239666 18226
rect 400 17782 239570 17894
rect 430 17778 239570 17782
rect 430 17666 239666 17778
rect 400 17446 239666 17666
rect 400 17330 239570 17446
rect 400 17222 239666 17330
rect 430 17106 239666 17222
rect 400 16998 239666 17106
rect 400 16882 239570 16998
rect 400 16662 239666 16882
rect 430 16550 239666 16662
rect 430 16546 239570 16550
rect 400 16434 239570 16546
rect 400 16102 239666 16434
rect 430 15986 239570 16102
rect 400 15654 239666 15986
rect 400 15542 239570 15654
rect 430 15538 239570 15542
rect 430 15426 239666 15538
rect 400 15206 239666 15426
rect 400 15090 239570 15206
rect 400 14982 239666 15090
rect 430 14866 239666 14982
rect 400 14758 239666 14866
rect 400 14642 239570 14758
rect 400 14422 239666 14642
rect 430 14310 239666 14422
rect 430 14306 239570 14310
rect 400 14194 239570 14306
rect 400 13862 239666 14194
rect 430 13746 239570 13862
rect 400 13414 239666 13746
rect 400 13302 239570 13414
rect 430 13298 239570 13302
rect 430 13186 239666 13298
rect 400 12966 239666 13186
rect 400 12850 239570 12966
rect 400 12742 239666 12850
rect 430 12626 239666 12742
rect 400 12518 239666 12626
rect 400 12402 239570 12518
rect 400 12182 239666 12402
rect 430 12070 239666 12182
rect 430 12066 239570 12070
rect 400 11954 239570 12066
rect 400 11622 239666 11954
rect 430 11506 239570 11622
rect 400 11174 239666 11506
rect 400 11062 239570 11174
rect 430 11058 239570 11062
rect 430 10946 239666 11058
rect 400 10726 239666 10946
rect 400 10610 239570 10726
rect 400 10502 239666 10610
rect 430 10386 239666 10502
rect 400 10278 239666 10386
rect 400 10162 239570 10278
rect 400 9942 239666 10162
rect 430 9830 239666 9942
rect 430 9826 239570 9830
rect 400 9714 239570 9826
rect 400 9382 239666 9714
rect 430 9266 239570 9382
rect 400 8934 239666 9266
rect 400 8822 239570 8934
rect 430 8818 239570 8822
rect 430 8706 239666 8818
rect 400 8486 239666 8706
rect 400 8370 239570 8486
rect 400 8262 239666 8370
rect 430 8146 239666 8262
rect 400 8038 239666 8146
rect 400 7922 239570 8038
rect 400 7702 239666 7922
rect 430 7590 239666 7702
rect 430 7586 239570 7590
rect 400 7474 239570 7586
rect 400 7142 239666 7474
rect 430 7026 239570 7142
rect 400 6694 239666 7026
rect 400 6582 239570 6694
rect 430 6578 239570 6582
rect 430 6466 239666 6578
rect 400 6246 239666 6466
rect 400 6130 239570 6246
rect 400 6022 239666 6130
rect 430 5906 239666 6022
rect 400 5798 239666 5906
rect 400 5682 239570 5798
rect 400 5462 239666 5682
rect 430 5350 239666 5462
rect 430 5346 239570 5350
rect 400 5234 239570 5346
rect 400 4902 239666 5234
rect 430 4786 239570 4902
rect 400 4454 239666 4786
rect 400 4342 239570 4454
rect 430 4338 239570 4342
rect 430 4226 239666 4338
rect 400 4006 239666 4226
rect 400 3890 239570 4006
rect 400 3782 239666 3890
rect 430 3666 239666 3782
rect 400 3558 239666 3666
rect 400 3442 239570 3558
rect 400 3222 239666 3442
rect 430 3110 239666 3222
rect 430 3106 239570 3110
rect 400 2994 239570 3106
rect 400 2662 239666 2994
rect 430 2546 239570 2662
rect 400 2214 239666 2546
rect 400 2102 239570 2214
rect 430 2098 239570 2102
rect 430 1986 239666 2098
rect 400 1766 239666 1986
rect 400 1650 239570 1766
rect 400 1318 239666 1650
rect 400 1202 239570 1318
rect 400 870 239666 1202
rect 400 754 239570 870
rect 400 238 239666 754
<< metal4 >>
rect 2224 1538 2384 28254
rect 9904 1538 10064 28254
rect 17584 1538 17744 28254
rect 25264 1538 25424 28254
rect 32944 1538 33104 28254
rect 40624 1538 40784 28254
rect 48304 1538 48464 28254
rect 55984 1538 56144 28254
rect 63664 1538 63824 28254
rect 71344 1538 71504 28254
rect 79024 1538 79184 28254
rect 86704 1538 86864 28254
rect 94384 1538 94544 28254
rect 102064 1538 102224 28254
rect 109744 1538 109904 28254
rect 117424 1538 117584 28254
rect 125104 1538 125264 28254
rect 132784 1538 132944 28254
rect 140464 1538 140624 28254
rect 148144 1538 148304 28254
rect 155824 1538 155984 28254
rect 163504 1538 163664 28254
rect 171184 1538 171344 28254
rect 178864 1538 179024 28254
rect 186544 1538 186704 28254
rect 194224 1538 194384 28254
rect 201904 1538 202064 28254
rect 209584 1538 209744 28254
rect 217264 1538 217424 28254
rect 224944 1538 225104 28254
rect 232624 1538 232784 28254
<< obsm4 >>
rect 69398 2081 71314 27711
rect 71534 2081 78994 27711
rect 79214 2081 86674 27711
rect 86894 2081 94354 27711
rect 94574 2081 102034 27711
rect 102254 2081 109714 27711
rect 109934 2081 117394 27711
rect 117614 2081 125074 27711
rect 125294 2081 132754 27711
rect 132974 2081 140434 27711
rect 140654 2081 148114 27711
rect 148334 2081 155794 27711
rect 156014 2081 163474 27711
rect 163694 2081 171154 27711
rect 171374 2081 172018 27711
<< labels >>
rlabel metal2 s 143472 0 143528 400 6 diego_clk
port 1 nsew signal output
rlabel metal2 s 144816 0 144872 400 6 diego_ena
port 2 nsew signal output
rlabel metal2 s 188496 0 188552 400 6 diego_io_in[0]
port 3 nsew signal output
rlabel metal2 s 195216 0 195272 400 6 diego_io_in[10]
port 4 nsew signal output
rlabel metal2 s 195888 0 195944 400 6 diego_io_in[11]
port 5 nsew signal output
rlabel metal2 s 196560 0 196616 400 6 diego_io_in[12]
port 6 nsew signal output
rlabel metal2 s 197232 0 197288 400 6 diego_io_in[13]
port 7 nsew signal output
rlabel metal2 s 197904 0 197960 400 6 diego_io_in[14]
port 8 nsew signal output
rlabel metal2 s 198576 0 198632 400 6 diego_io_in[15]
port 9 nsew signal output
rlabel metal2 s 199248 0 199304 400 6 diego_io_in[16]
port 10 nsew signal output
rlabel metal2 s 199920 0 199976 400 6 diego_io_in[17]
port 11 nsew signal output
rlabel metal2 s 200592 0 200648 400 6 diego_io_in[18]
port 12 nsew signal output
rlabel metal2 s 201264 0 201320 400 6 diego_io_in[19]
port 13 nsew signal output
rlabel metal2 s 189168 0 189224 400 6 diego_io_in[1]
port 14 nsew signal output
rlabel metal2 s 201936 0 201992 400 6 diego_io_in[20]
port 15 nsew signal output
rlabel metal2 s 202608 0 202664 400 6 diego_io_in[21]
port 16 nsew signal output
rlabel metal2 s 203280 0 203336 400 6 diego_io_in[22]
port 17 nsew signal output
rlabel metal2 s 203952 0 204008 400 6 diego_io_in[23]
port 18 nsew signal output
rlabel metal2 s 204624 0 204680 400 6 diego_io_in[24]
port 19 nsew signal output
rlabel metal2 s 205296 0 205352 400 6 diego_io_in[25]
port 20 nsew signal output
rlabel metal2 s 205968 0 206024 400 6 diego_io_in[26]
port 21 nsew signal output
rlabel metal2 s 206640 0 206696 400 6 diego_io_in[27]
port 22 nsew signal output
rlabel metal2 s 207312 0 207368 400 6 diego_io_in[28]
port 23 nsew signal output
rlabel metal2 s 207984 0 208040 400 6 diego_io_in[29]
port 24 nsew signal output
rlabel metal2 s 189840 0 189896 400 6 diego_io_in[2]
port 25 nsew signal output
rlabel metal2 s 208656 0 208712 400 6 diego_io_in[30]
port 26 nsew signal output
rlabel metal2 s 209328 0 209384 400 6 diego_io_in[31]
port 27 nsew signal output
rlabel metal2 s 210000 0 210056 400 6 diego_io_in[32]
port 28 nsew signal output
rlabel metal2 s 210672 0 210728 400 6 diego_io_in[33]
port 29 nsew signal output
rlabel metal2 s 211344 0 211400 400 6 diego_io_in[34]
port 30 nsew signal output
rlabel metal2 s 212016 0 212072 400 6 diego_io_in[35]
port 31 nsew signal output
rlabel metal2 s 212688 0 212744 400 6 diego_io_in[36]
port 32 nsew signal output
rlabel metal2 s 213360 0 213416 400 6 diego_io_in[37]
port 33 nsew signal output
rlabel metal2 s 190512 0 190568 400 6 diego_io_in[3]
port 34 nsew signal output
rlabel metal2 s 191184 0 191240 400 6 diego_io_in[4]
port 35 nsew signal output
rlabel metal2 s 191856 0 191912 400 6 diego_io_in[5]
port 36 nsew signal output
rlabel metal2 s 192528 0 192584 400 6 diego_io_in[6]
port 37 nsew signal output
rlabel metal2 s 193200 0 193256 400 6 diego_io_in[7]
port 38 nsew signal output
rlabel metal2 s 193872 0 193928 400 6 diego_io_in[8]
port 39 nsew signal output
rlabel metal2 s 194544 0 194600 400 6 diego_io_in[9]
port 40 nsew signal output
rlabel metal2 s 166992 0 167048 400 6 diego_io_oeb[0]
port 41 nsew signal input
rlabel metal2 s 173712 0 173768 400 6 diego_io_oeb[10]
port 42 nsew signal input
rlabel metal2 s 174384 0 174440 400 6 diego_io_oeb[11]
port 43 nsew signal input
rlabel metal2 s 175056 0 175112 400 6 diego_io_oeb[12]
port 44 nsew signal input
rlabel metal2 s 175728 0 175784 400 6 diego_io_oeb[13]
port 45 nsew signal input
rlabel metal2 s 176400 0 176456 400 6 diego_io_oeb[14]
port 46 nsew signal input
rlabel metal2 s 177072 0 177128 400 6 diego_io_oeb[15]
port 47 nsew signal input
rlabel metal2 s 177744 0 177800 400 6 diego_io_oeb[16]
port 48 nsew signal input
rlabel metal2 s 178416 0 178472 400 6 diego_io_oeb[17]
port 49 nsew signal input
rlabel metal2 s 179088 0 179144 400 6 diego_io_oeb[18]
port 50 nsew signal input
rlabel metal2 s 179760 0 179816 400 6 diego_io_oeb[19]
port 51 nsew signal input
rlabel metal2 s 167664 0 167720 400 6 diego_io_oeb[1]
port 52 nsew signal input
rlabel metal2 s 180432 0 180488 400 6 diego_io_oeb[20]
port 53 nsew signal input
rlabel metal2 s 181104 0 181160 400 6 diego_io_oeb[21]
port 54 nsew signal input
rlabel metal2 s 181776 0 181832 400 6 diego_io_oeb[22]
port 55 nsew signal input
rlabel metal2 s 182448 0 182504 400 6 diego_io_oeb[23]
port 56 nsew signal input
rlabel metal2 s 183120 0 183176 400 6 diego_io_oeb[24]
port 57 nsew signal input
rlabel metal2 s 183792 0 183848 400 6 diego_io_oeb[25]
port 58 nsew signal input
rlabel metal2 s 184464 0 184520 400 6 diego_io_oeb[26]
port 59 nsew signal input
rlabel metal2 s 185136 0 185192 400 6 diego_io_oeb[27]
port 60 nsew signal input
rlabel metal2 s 185808 0 185864 400 6 diego_io_oeb[28]
port 61 nsew signal input
rlabel metal2 s 186480 0 186536 400 6 diego_io_oeb[29]
port 62 nsew signal input
rlabel metal2 s 168336 0 168392 400 6 diego_io_oeb[2]
port 63 nsew signal input
rlabel metal2 s 187152 0 187208 400 6 diego_io_oeb[30]
port 64 nsew signal input
rlabel metal2 s 187824 0 187880 400 6 diego_io_oeb[31]
port 65 nsew signal input
rlabel metal2 s 169008 0 169064 400 6 diego_io_oeb[3]
port 66 nsew signal input
rlabel metal2 s 169680 0 169736 400 6 diego_io_oeb[4]
port 67 nsew signal input
rlabel metal2 s 170352 0 170408 400 6 diego_io_oeb[5]
port 68 nsew signal input
rlabel metal2 s 171024 0 171080 400 6 diego_io_oeb[6]
port 69 nsew signal input
rlabel metal2 s 171696 0 171752 400 6 diego_io_oeb[7]
port 70 nsew signal input
rlabel metal2 s 172368 0 172424 400 6 diego_io_oeb[8]
port 71 nsew signal input
rlabel metal2 s 173040 0 173096 400 6 diego_io_oeb[9]
port 72 nsew signal input
rlabel metal2 s 145488 0 145544 400 6 diego_io_out[0]
port 73 nsew signal input
rlabel metal2 s 152208 0 152264 400 6 diego_io_out[10]
port 74 nsew signal input
rlabel metal2 s 152880 0 152936 400 6 diego_io_out[11]
port 75 nsew signal input
rlabel metal2 s 153552 0 153608 400 6 diego_io_out[12]
port 76 nsew signal input
rlabel metal2 s 154224 0 154280 400 6 diego_io_out[13]
port 77 nsew signal input
rlabel metal2 s 154896 0 154952 400 6 diego_io_out[14]
port 78 nsew signal input
rlabel metal2 s 155568 0 155624 400 6 diego_io_out[15]
port 79 nsew signal input
rlabel metal2 s 156240 0 156296 400 6 diego_io_out[16]
port 80 nsew signal input
rlabel metal2 s 156912 0 156968 400 6 diego_io_out[17]
port 81 nsew signal input
rlabel metal2 s 157584 0 157640 400 6 diego_io_out[18]
port 82 nsew signal input
rlabel metal2 s 158256 0 158312 400 6 diego_io_out[19]
port 83 nsew signal input
rlabel metal2 s 146160 0 146216 400 6 diego_io_out[1]
port 84 nsew signal input
rlabel metal2 s 158928 0 158984 400 6 diego_io_out[20]
port 85 nsew signal input
rlabel metal2 s 159600 0 159656 400 6 diego_io_out[21]
port 86 nsew signal input
rlabel metal2 s 160272 0 160328 400 6 diego_io_out[22]
port 87 nsew signal input
rlabel metal2 s 160944 0 161000 400 6 diego_io_out[23]
port 88 nsew signal input
rlabel metal2 s 161616 0 161672 400 6 diego_io_out[24]
port 89 nsew signal input
rlabel metal2 s 162288 0 162344 400 6 diego_io_out[25]
port 90 nsew signal input
rlabel metal2 s 162960 0 163016 400 6 diego_io_out[26]
port 91 nsew signal input
rlabel metal2 s 163632 0 163688 400 6 diego_io_out[27]
port 92 nsew signal input
rlabel metal2 s 164304 0 164360 400 6 diego_io_out[28]
port 93 nsew signal input
rlabel metal2 s 164976 0 165032 400 6 diego_io_out[29]
port 94 nsew signal input
rlabel metal2 s 146832 0 146888 400 6 diego_io_out[2]
port 95 nsew signal input
rlabel metal2 s 165648 0 165704 400 6 diego_io_out[30]
port 96 nsew signal input
rlabel metal2 s 166320 0 166376 400 6 diego_io_out[31]
port 97 nsew signal input
rlabel metal2 s 147504 0 147560 400 6 diego_io_out[3]
port 98 nsew signal input
rlabel metal2 s 148176 0 148232 400 6 diego_io_out[4]
port 99 nsew signal input
rlabel metal2 s 148848 0 148904 400 6 diego_io_out[5]
port 100 nsew signal input
rlabel metal2 s 149520 0 149576 400 6 diego_io_out[6]
port 101 nsew signal input
rlabel metal2 s 150192 0 150248 400 6 diego_io_out[7]
port 102 nsew signal input
rlabel metal2 s 150864 0 150920 400 6 diego_io_out[8]
port 103 nsew signal input
rlabel metal2 s 151536 0 151592 400 6 diego_io_out[9]
port 104 nsew signal input
rlabel metal2 s 144144 0 144200 400 6 diego_rst
port 105 nsew signal output
rlabel metal3 s 239600 3920 240000 3976 6 i_design_reset[0]
port 106 nsew signal input
rlabel metal3 s 239600 4368 240000 4424 6 i_design_reset[1]
port 107 nsew signal input
rlabel metal3 s 239600 4816 240000 4872 6 i_design_reset[2]
port 108 nsew signal input
rlabel metal3 s 239600 5264 240000 5320 6 i_design_reset[3]
port 109 nsew signal input
rlabel metal3 s 239600 5712 240000 5768 6 i_design_reset[4]
port 110 nsew signal input
rlabel metal3 s 239600 6160 240000 6216 6 i_design_reset[5]
port 111 nsew signal input
rlabel metal3 s 239600 6608 240000 6664 6 i_design_reset[6]
port 112 nsew signal input
rlabel metal3 s 239600 7056 240000 7112 6 i_design_reset[7]
port 113 nsew signal input
rlabel metal3 s 239600 3472 240000 3528 6 i_mux_auto_reset_enb
port 114 nsew signal input
rlabel metal3 s 239600 784 240000 840 6 i_mux_io5_reset_enb
port 115 nsew signal input
rlabel metal3 s 239600 1232 240000 1288 6 i_mux_sel[0]
port 116 nsew signal input
rlabel metal3 s 239600 1680 240000 1736 6 i_mux_sel[1]
port 117 nsew signal input
rlabel metal3 s 239600 2128 240000 2184 6 i_mux_sel[2]
port 118 nsew signal input
rlabel metal3 s 239600 2576 240000 2632 6 i_mux_sel[3]
port 119 nsew signal input
rlabel metal3 s 239600 3024 240000 3080 6 i_mux_sys_reset_enb
port 120 nsew signal input
rlabel metal3 s 239600 7952 240000 8008 6 io_in[0]
port 121 nsew signal input
rlabel metal3 s 239600 21392 240000 21448 6 io_in[10]
port 122 nsew signal input
rlabel metal3 s 239600 22736 240000 22792 6 io_in[11]
port 123 nsew signal input
rlabel metal3 s 239600 24080 240000 24136 6 io_in[12]
port 124 nsew signal input
rlabel metal3 s 239600 25424 240000 25480 6 io_in[13]
port 125 nsew signal input
rlabel metal3 s 239600 26768 240000 26824 6 io_in[14]
port 126 nsew signal input
rlabel metal3 s 239600 28112 240000 28168 6 io_in[15]
port 127 nsew signal input
rlabel metal2 s 196224 29600 196280 30000 6 io_in[16]
port 128 nsew signal input
rlabel metal2 s 194208 29600 194264 30000 6 io_in[17]
port 129 nsew signal input
rlabel metal2 s 192192 29600 192248 30000 6 io_in[18]
port 130 nsew signal input
rlabel metal2 s 63840 29600 63896 30000 6 io_in[19]
port 131 nsew signal input
rlabel metal3 s 239600 9296 240000 9352 6 io_in[1]
port 132 nsew signal input
rlabel metal2 s 61824 29600 61880 30000 6 io_in[20]
port 133 nsew signal input
rlabel metal2 s 59808 29600 59864 30000 6 io_in[21]
port 134 nsew signal input
rlabel metal2 s 57792 29600 57848 30000 6 io_in[22]
port 135 nsew signal input
rlabel metal3 s 0 27776 400 27832 6 io_in[23]
port 136 nsew signal input
rlabel metal3 s 0 26096 400 26152 6 io_in[24]
port 137 nsew signal input
rlabel metal3 s 0 24416 400 24472 6 io_in[25]
port 138 nsew signal input
rlabel metal3 s 0 22736 400 22792 6 io_in[26]
port 139 nsew signal input
rlabel metal3 s 0 21056 400 21112 6 io_in[27]
port 140 nsew signal input
rlabel metal3 s 0 19376 400 19432 6 io_in[28]
port 141 nsew signal input
rlabel metal3 s 0 17696 400 17752 6 io_in[29]
port 142 nsew signal input
rlabel metal3 s 239600 10640 240000 10696 6 io_in[2]
port 143 nsew signal input
rlabel metal3 s 0 16016 400 16072 6 io_in[30]
port 144 nsew signal input
rlabel metal3 s 0 14336 400 14392 6 io_in[31]
port 145 nsew signal input
rlabel metal3 s 0 12656 400 12712 6 io_in[32]
port 146 nsew signal input
rlabel metal3 s 0 10976 400 11032 6 io_in[33]
port 147 nsew signal input
rlabel metal3 s 0 9296 400 9352 6 io_in[34]
port 148 nsew signal input
rlabel metal3 s 0 7616 400 7672 6 io_in[35]
port 149 nsew signal input
rlabel metal3 s 0 5936 400 5992 6 io_in[36]
port 150 nsew signal input
rlabel metal3 s 0 4256 400 4312 6 io_in[37]
port 151 nsew signal input
rlabel metal3 s 239600 11984 240000 12040 6 io_in[3]
port 152 nsew signal input
rlabel metal3 s 239600 13328 240000 13384 6 io_in[4]
port 153 nsew signal input
rlabel metal3 s 239600 14672 240000 14728 6 io_in[5]
port 154 nsew signal input
rlabel metal3 s 239600 16016 240000 16072 6 io_in[6]
port 155 nsew signal input
rlabel metal3 s 239600 17360 240000 17416 6 io_in[7]
port 156 nsew signal input
rlabel metal3 s 239600 18704 240000 18760 6 io_in[8]
port 157 nsew signal input
rlabel metal3 s 239600 20048 240000 20104 6 io_in[9]
port 158 nsew signal input
rlabel metal3 s 239600 8848 240000 8904 6 io_oeb[0]
port 159 nsew signal output
rlabel metal3 s 239600 22288 240000 22344 6 io_oeb[10]
port 160 nsew signal output
rlabel metal3 s 239600 23632 240000 23688 6 io_oeb[11]
port 161 nsew signal output
rlabel metal3 s 239600 24976 240000 25032 6 io_oeb[12]
port 162 nsew signal output
rlabel metal3 s 239600 26320 240000 26376 6 io_oeb[13]
port 163 nsew signal output
rlabel metal3 s 239600 27664 240000 27720 6 io_oeb[14]
port 164 nsew signal output
rlabel metal3 s 239600 29008 240000 29064 6 io_oeb[15]
port 165 nsew signal output
rlabel metal2 s 194880 29600 194936 30000 6 io_oeb[16]
port 166 nsew signal output
rlabel metal2 s 192864 29600 192920 30000 6 io_oeb[17]
port 167 nsew signal output
rlabel metal2 s 190848 29600 190904 30000 6 io_oeb[18]
port 168 nsew signal output
rlabel metal2 s 62496 29600 62552 30000 6 io_oeb[19]
port 169 nsew signal output
rlabel metal3 s 239600 10192 240000 10248 6 io_oeb[1]
port 170 nsew signal output
rlabel metal2 s 60480 29600 60536 30000 6 io_oeb[20]
port 171 nsew signal output
rlabel metal2 s 58464 29600 58520 30000 6 io_oeb[21]
port 172 nsew signal output
rlabel metal2 s 56448 29600 56504 30000 6 io_oeb[22]
port 173 nsew signal output
rlabel metal3 s 0 26656 400 26712 6 io_oeb[23]
port 174 nsew signal output
rlabel metal3 s 0 24976 400 25032 6 io_oeb[24]
port 175 nsew signal output
rlabel metal3 s 0 23296 400 23352 6 io_oeb[25]
port 176 nsew signal output
rlabel metal3 s 0 21616 400 21672 6 io_oeb[26]
port 177 nsew signal output
rlabel metal3 s 0 19936 400 19992 6 io_oeb[27]
port 178 nsew signal output
rlabel metal3 s 0 18256 400 18312 6 io_oeb[28]
port 179 nsew signal output
rlabel metal3 s 0 16576 400 16632 6 io_oeb[29]
port 180 nsew signal output
rlabel metal3 s 239600 11536 240000 11592 6 io_oeb[2]
port 181 nsew signal output
rlabel metal3 s 0 14896 400 14952 6 io_oeb[30]
port 182 nsew signal output
rlabel metal3 s 0 13216 400 13272 6 io_oeb[31]
port 183 nsew signal output
rlabel metal3 s 0 11536 400 11592 6 io_oeb[32]
port 184 nsew signal output
rlabel metal3 s 0 9856 400 9912 6 io_oeb[33]
port 185 nsew signal output
rlabel metal3 s 0 8176 400 8232 6 io_oeb[34]
port 186 nsew signal output
rlabel metal3 s 0 6496 400 6552 6 io_oeb[35]
port 187 nsew signal output
rlabel metal3 s 0 4816 400 4872 6 io_oeb[36]
port 188 nsew signal output
rlabel metal3 s 0 3136 400 3192 6 io_oeb[37]
port 189 nsew signal output
rlabel metal3 s 239600 12880 240000 12936 6 io_oeb[3]
port 190 nsew signal output
rlabel metal3 s 239600 14224 240000 14280 6 io_oeb[4]
port 191 nsew signal output
rlabel metal3 s 239600 15568 240000 15624 6 io_oeb[5]
port 192 nsew signal output
rlabel metal3 s 239600 16912 240000 16968 6 io_oeb[6]
port 193 nsew signal output
rlabel metal3 s 239600 18256 240000 18312 6 io_oeb[7]
port 194 nsew signal output
rlabel metal3 s 239600 19600 240000 19656 6 io_oeb[8]
port 195 nsew signal output
rlabel metal3 s 239600 20944 240000 21000 6 io_oeb[9]
port 196 nsew signal output
rlabel metal3 s 239600 8400 240000 8456 6 io_out[0]
port 197 nsew signal output
rlabel metal3 s 239600 21840 240000 21896 6 io_out[10]
port 198 nsew signal output
rlabel metal3 s 239600 23184 240000 23240 6 io_out[11]
port 199 nsew signal output
rlabel metal3 s 239600 24528 240000 24584 6 io_out[12]
port 200 nsew signal output
rlabel metal3 s 239600 25872 240000 25928 6 io_out[13]
port 201 nsew signal output
rlabel metal3 s 239600 27216 240000 27272 6 io_out[14]
port 202 nsew signal output
rlabel metal3 s 239600 28560 240000 28616 6 io_out[15]
port 203 nsew signal output
rlabel metal2 s 195552 29600 195608 30000 6 io_out[16]
port 204 nsew signal output
rlabel metal2 s 193536 29600 193592 30000 6 io_out[17]
port 205 nsew signal output
rlabel metal2 s 191520 29600 191576 30000 6 io_out[18]
port 206 nsew signal output
rlabel metal2 s 63168 29600 63224 30000 6 io_out[19]
port 207 nsew signal output
rlabel metal3 s 239600 9744 240000 9800 6 io_out[1]
port 208 nsew signal output
rlabel metal2 s 61152 29600 61208 30000 6 io_out[20]
port 209 nsew signal output
rlabel metal2 s 59136 29600 59192 30000 6 io_out[21]
port 210 nsew signal output
rlabel metal2 s 57120 29600 57176 30000 6 io_out[22]
port 211 nsew signal output
rlabel metal3 s 0 27216 400 27272 6 io_out[23]
port 212 nsew signal output
rlabel metal3 s 0 25536 400 25592 6 io_out[24]
port 213 nsew signal output
rlabel metal3 s 0 23856 400 23912 6 io_out[25]
port 214 nsew signal output
rlabel metal3 s 0 22176 400 22232 6 io_out[26]
port 215 nsew signal output
rlabel metal3 s 0 20496 400 20552 6 io_out[27]
port 216 nsew signal output
rlabel metal3 s 0 18816 400 18872 6 io_out[28]
port 217 nsew signal output
rlabel metal3 s 0 17136 400 17192 6 io_out[29]
port 218 nsew signal output
rlabel metal3 s 239600 11088 240000 11144 6 io_out[2]
port 219 nsew signal output
rlabel metal3 s 0 15456 400 15512 6 io_out[30]
port 220 nsew signal output
rlabel metal3 s 0 13776 400 13832 6 io_out[31]
port 221 nsew signal output
rlabel metal3 s 0 12096 400 12152 6 io_out[32]
port 222 nsew signal output
rlabel metal3 s 0 10416 400 10472 6 io_out[33]
port 223 nsew signal output
rlabel metal3 s 0 8736 400 8792 6 io_out[34]
port 224 nsew signal output
rlabel metal3 s 0 7056 400 7112 6 io_out[35]
port 225 nsew signal output
rlabel metal3 s 0 5376 400 5432 6 io_out[36]
port 226 nsew signal output
rlabel metal3 s 0 3696 400 3752 6 io_out[37]
port 227 nsew signal output
rlabel metal3 s 239600 12432 240000 12488 6 io_out[3]
port 228 nsew signal output
rlabel metal3 s 239600 13776 240000 13832 6 io_out[4]
port 229 nsew signal output
rlabel metal3 s 239600 15120 240000 15176 6 io_out[5]
port 230 nsew signal output
rlabel metal3 s 239600 16464 240000 16520 6 io_out[6]
port 231 nsew signal output
rlabel metal3 s 239600 17808 240000 17864 6 io_out[7]
port 232 nsew signal output
rlabel metal3 s 239600 19152 240000 19208 6 io_out[8]
port 233 nsew signal output
rlabel metal3 s 239600 20496 240000 20552 6 io_out[9]
port 234 nsew signal output
rlabel metal2 s 112560 0 112616 400 6 la_in[0]
port 235 nsew signal input
rlabel metal2 s 119280 0 119336 400 6 la_in[10]
port 236 nsew signal input
rlabel metal2 s 119952 0 120008 400 6 la_in[11]
port 237 nsew signal input
rlabel metal2 s 120624 0 120680 400 6 la_in[12]
port 238 nsew signal input
rlabel metal2 s 121296 0 121352 400 6 la_in[13]
port 239 nsew signal input
rlabel metal2 s 121968 0 122024 400 6 la_in[14]
port 240 nsew signal input
rlabel metal2 s 122640 0 122696 400 6 la_in[15]
port 241 nsew signal input
rlabel metal2 s 113232 0 113288 400 6 la_in[1]
port 242 nsew signal input
rlabel metal2 s 113904 0 113960 400 6 la_in[2]
port 243 nsew signal input
rlabel metal2 s 114576 0 114632 400 6 la_in[3]
port 244 nsew signal input
rlabel metal2 s 115248 0 115304 400 6 la_in[4]
port 245 nsew signal input
rlabel metal2 s 115920 0 115976 400 6 la_in[5]
port 246 nsew signal input
rlabel metal2 s 116592 0 116648 400 6 la_in[6]
port 247 nsew signal input
rlabel metal2 s 117264 0 117320 400 6 la_in[7]
port 248 nsew signal input
rlabel metal2 s 117936 0 117992 400 6 la_in[8]
port 249 nsew signal input
rlabel metal2 s 118608 0 118664 400 6 la_in[9]
port 250 nsew signal input
rlabel metal3 s 239600 7504 240000 7560 6 mux_conf_clk
port 251 nsew signal input
rlabel metal2 s 4368 0 4424 400 6 pawel_clk
port 252 nsew signal output
rlabel metal2 s 5712 0 5768 400 6 pawel_ena
port 253 nsew signal output
rlabel metal2 s 6384 0 6440 400 6 pawel_io_in[0]
port 254 nsew signal output
rlabel metal2 s 26544 0 26600 400 6 pawel_io_in[10]
port 255 nsew signal output
rlabel metal2 s 28560 0 28616 400 6 pawel_io_in[11]
port 256 nsew signal output
rlabel metal2 s 30576 0 30632 400 6 pawel_io_in[12]
port 257 nsew signal output
rlabel metal2 s 32592 0 32648 400 6 pawel_io_in[13]
port 258 nsew signal output
rlabel metal2 s 33264 0 33320 400 6 pawel_io_in[14]
port 259 nsew signal output
rlabel metal2 s 33936 0 33992 400 6 pawel_io_in[15]
port 260 nsew signal output
rlabel metal2 s 34608 0 34664 400 6 pawel_io_in[16]
port 261 nsew signal output
rlabel metal2 s 35280 0 35336 400 6 pawel_io_in[17]
port 262 nsew signal output
rlabel metal2 s 35952 0 36008 400 6 pawel_io_in[18]
port 263 nsew signal output
rlabel metal2 s 36624 0 36680 400 6 pawel_io_in[19]
port 264 nsew signal output
rlabel metal2 s 8400 0 8456 400 6 pawel_io_in[1]
port 265 nsew signal output
rlabel metal2 s 37296 0 37352 400 6 pawel_io_in[20]
port 266 nsew signal output
rlabel metal2 s 37968 0 38024 400 6 pawel_io_in[21]
port 267 nsew signal output
rlabel metal2 s 38640 0 38696 400 6 pawel_io_in[22]
port 268 nsew signal output
rlabel metal2 s 39312 0 39368 400 6 pawel_io_in[23]
port 269 nsew signal output
rlabel metal2 s 39984 0 40040 400 6 pawel_io_in[24]
port 270 nsew signal output
rlabel metal2 s 40656 0 40712 400 6 pawel_io_in[25]
port 271 nsew signal output
rlabel metal2 s 41328 0 41384 400 6 pawel_io_in[26]
port 272 nsew signal output
rlabel metal2 s 42000 0 42056 400 6 pawel_io_in[27]
port 273 nsew signal output
rlabel metal2 s 42672 0 42728 400 6 pawel_io_in[28]
port 274 nsew signal output
rlabel metal2 s 43344 0 43400 400 6 pawel_io_in[29]
port 275 nsew signal output
rlabel metal2 s 10416 0 10472 400 6 pawel_io_in[2]
port 276 nsew signal output
rlabel metal2 s 44016 0 44072 400 6 pawel_io_in[30]
port 277 nsew signal output
rlabel metal2 s 44688 0 44744 400 6 pawel_io_in[31]
port 278 nsew signal output
rlabel metal2 s 45360 0 45416 400 6 pawel_io_in[32]
port 279 nsew signal output
rlabel metal2 s 46032 0 46088 400 6 pawel_io_in[33]
port 280 nsew signal output
rlabel metal2 s 46704 0 46760 400 6 pawel_io_in[34]
port 281 nsew signal output
rlabel metal2 s 47376 0 47432 400 6 pawel_io_in[35]
port 282 nsew signal output
rlabel metal2 s 48048 0 48104 400 6 pawel_io_in[36]
port 283 nsew signal output
rlabel metal2 s 48720 0 48776 400 6 pawel_io_in[37]
port 284 nsew signal output
rlabel metal2 s 12432 0 12488 400 6 pawel_io_in[3]
port 285 nsew signal output
rlabel metal2 s 14448 0 14504 400 6 pawel_io_in[4]
port 286 nsew signal output
rlabel metal2 s 16464 0 16520 400 6 pawel_io_in[5]
port 287 nsew signal output
rlabel metal2 s 18480 0 18536 400 6 pawel_io_in[6]
port 288 nsew signal output
rlabel metal2 s 20496 0 20552 400 6 pawel_io_in[7]
port 289 nsew signal output
rlabel metal2 s 22512 0 22568 400 6 pawel_io_in[8]
port 290 nsew signal output
rlabel metal2 s 24528 0 24584 400 6 pawel_io_in[9]
port 291 nsew signal output
rlabel metal2 s 7056 0 7112 400 6 pawel_io_oeb[0]
port 292 nsew signal input
rlabel metal2 s 27216 0 27272 400 6 pawel_io_oeb[10]
port 293 nsew signal input
rlabel metal2 s 29232 0 29288 400 6 pawel_io_oeb[11]
port 294 nsew signal input
rlabel metal2 s 31248 0 31304 400 6 pawel_io_oeb[12]
port 295 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 pawel_io_oeb[1]
port 296 nsew signal input
rlabel metal2 s 11088 0 11144 400 6 pawel_io_oeb[2]
port 297 nsew signal input
rlabel metal2 s 13104 0 13160 400 6 pawel_io_oeb[3]
port 298 nsew signal input
rlabel metal2 s 15120 0 15176 400 6 pawel_io_oeb[4]
port 299 nsew signal input
rlabel metal2 s 17136 0 17192 400 6 pawel_io_oeb[5]
port 300 nsew signal input
rlabel metal2 s 19152 0 19208 400 6 pawel_io_oeb[6]
port 301 nsew signal input
rlabel metal2 s 21168 0 21224 400 6 pawel_io_oeb[7]
port 302 nsew signal input
rlabel metal2 s 23184 0 23240 400 6 pawel_io_oeb[8]
port 303 nsew signal input
rlabel metal2 s 25200 0 25256 400 6 pawel_io_oeb[9]
port 304 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 pawel_io_out[0]
port 305 nsew signal input
rlabel metal2 s 27888 0 27944 400 6 pawel_io_out[10]
port 306 nsew signal input
rlabel metal2 s 29904 0 29960 400 6 pawel_io_out[11]
port 307 nsew signal input
rlabel metal2 s 31920 0 31976 400 6 pawel_io_out[12]
port 308 nsew signal input
rlabel metal2 s 9744 0 9800 400 6 pawel_io_out[1]
port 309 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 pawel_io_out[2]
port 310 nsew signal input
rlabel metal2 s 13776 0 13832 400 6 pawel_io_out[3]
port 311 nsew signal input
rlabel metal2 s 15792 0 15848 400 6 pawel_io_out[4]
port 312 nsew signal input
rlabel metal2 s 17808 0 17864 400 6 pawel_io_out[5]
port 313 nsew signal input
rlabel metal2 s 19824 0 19880 400 6 pawel_io_out[6]
port 314 nsew signal input
rlabel metal2 s 21840 0 21896 400 6 pawel_io_out[7]
port 315 nsew signal input
rlabel metal2 s 23856 0 23912 400 6 pawel_io_out[8]
port 316 nsew signal input
rlabel metal2 s 25872 0 25928 400 6 pawel_io_out[9]
port 317 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 pawel_rst
port 318 nsew signal output
rlabel metal2 s 200256 29600 200312 30000 6 solos_clk
port 319 nsew signal output
rlabel metal2 s 201600 29600 201656 30000 6 solos_ena
port 320 nsew signal output
rlabel metal2 s 202272 29600 202328 30000 6 solos_gpio_ready
port 321 nsew signal output
rlabel metal2 s 236544 29600 236600 30000 6 solos_io_in[0]
port 322 nsew signal output
rlabel metal2 s 229824 29600 229880 30000 6 solos_io_in[10]
port 323 nsew signal output
rlabel metal2 s 229152 29600 229208 30000 6 solos_io_in[11]
port 324 nsew signal output
rlabel metal2 s 228480 29600 228536 30000 6 solos_io_in[12]
port 325 nsew signal output
rlabel metal2 s 227808 29600 227864 30000 6 solos_io_in[13]
port 326 nsew signal output
rlabel metal2 s 227136 29600 227192 30000 6 solos_io_in[14]
port 327 nsew signal output
rlabel metal2 s 226464 29600 226520 30000 6 solos_io_in[15]
port 328 nsew signal output
rlabel metal2 s 225792 29600 225848 30000 6 solos_io_in[16]
port 329 nsew signal output
rlabel metal2 s 225120 29600 225176 30000 6 solos_io_in[17]
port 330 nsew signal output
rlabel metal2 s 224448 29600 224504 30000 6 solos_io_in[18]
port 331 nsew signal output
rlabel metal2 s 223776 29600 223832 30000 6 solos_io_in[19]
port 332 nsew signal output
rlabel metal2 s 235872 29600 235928 30000 6 solos_io_in[1]
port 333 nsew signal output
rlabel metal2 s 223104 29600 223160 30000 6 solos_io_in[20]
port 334 nsew signal output
rlabel metal2 s 222432 29600 222488 30000 6 solos_io_in[21]
port 335 nsew signal output
rlabel metal2 s 221760 29600 221816 30000 6 solos_io_in[22]
port 336 nsew signal output
rlabel metal2 s 221088 29600 221144 30000 6 solos_io_in[23]
port 337 nsew signal output
rlabel metal2 s 220416 29600 220472 30000 6 solos_io_in[24]
port 338 nsew signal output
rlabel metal2 s 219744 29600 219800 30000 6 solos_io_in[25]
port 339 nsew signal output
rlabel metal2 s 219072 29600 219128 30000 6 solos_io_in[26]
port 340 nsew signal output
rlabel metal2 s 218400 29600 218456 30000 6 solos_io_in[27]
port 341 nsew signal output
rlabel metal2 s 217728 29600 217784 30000 6 solos_io_in[28]
port 342 nsew signal output
rlabel metal2 s 217056 29600 217112 30000 6 solos_io_in[29]
port 343 nsew signal output
rlabel metal2 s 235200 29600 235256 30000 6 solos_io_in[2]
port 344 nsew signal output
rlabel metal2 s 216384 29600 216440 30000 6 solos_io_in[30]
port 345 nsew signal output
rlabel metal2 s 215712 29600 215768 30000 6 solos_io_in[31]
port 346 nsew signal output
rlabel metal2 s 215040 29600 215096 30000 6 solos_io_in[32]
port 347 nsew signal output
rlabel metal2 s 214368 29600 214424 30000 6 solos_io_in[33]
port 348 nsew signal output
rlabel metal2 s 213696 29600 213752 30000 6 solos_io_in[34]
port 349 nsew signal output
rlabel metal2 s 213024 29600 213080 30000 6 solos_io_in[35]
port 350 nsew signal output
rlabel metal2 s 212352 29600 212408 30000 6 solos_io_in[36]
port 351 nsew signal output
rlabel metal2 s 211680 29600 211736 30000 6 solos_io_in[37]
port 352 nsew signal output
rlabel metal2 s 234528 29600 234584 30000 6 solos_io_in[3]
port 353 nsew signal output
rlabel metal2 s 233856 29600 233912 30000 6 solos_io_in[4]
port 354 nsew signal output
rlabel metal2 s 233184 29600 233240 30000 6 solos_io_in[5]
port 355 nsew signal output
rlabel metal2 s 232512 29600 232568 30000 6 solos_io_in[6]
port 356 nsew signal output
rlabel metal2 s 231840 29600 231896 30000 6 solos_io_in[7]
port 357 nsew signal output
rlabel metal2 s 231168 29600 231224 30000 6 solos_io_in[8]
port 358 nsew signal output
rlabel metal2 s 230496 29600 230552 30000 6 solos_io_in[9]
port 359 nsew signal output
rlabel metal2 s 211008 29600 211064 30000 6 solos_io_out[0]
port 360 nsew signal input
rlabel metal2 s 204288 29600 204344 30000 6 solos_io_out[10]
port 361 nsew signal input
rlabel metal2 s 203616 29600 203672 30000 6 solos_io_out[11]
port 362 nsew signal input
rlabel metal2 s 202944 29600 203000 30000 6 solos_io_out[12]
port 363 nsew signal input
rlabel metal2 s 210336 29600 210392 30000 6 solos_io_out[1]
port 364 nsew signal input
rlabel metal2 s 209664 29600 209720 30000 6 solos_io_out[2]
port 365 nsew signal input
rlabel metal2 s 208992 29600 209048 30000 6 solos_io_out[3]
port 366 nsew signal input
rlabel metal2 s 208320 29600 208376 30000 6 solos_io_out[4]
port 367 nsew signal input
rlabel metal2 s 207648 29600 207704 30000 6 solos_io_out[5]
port 368 nsew signal input
rlabel metal2 s 206976 29600 207032 30000 6 solos_io_out[6]
port 369 nsew signal input
rlabel metal2 s 206304 29600 206360 30000 6 solos_io_out[7]
port 370 nsew signal input
rlabel metal2 s 205632 29600 205688 30000 6 solos_io_out[8]
port 371 nsew signal input
rlabel metal2 s 204960 29600 205016 30000 6 solos_io_out[9]
port 372 nsew signal input
rlabel metal2 s 200928 29600 200984 30000 6 solos_rst
port 373 nsew signal output
rlabel metal2 s 71904 29600 71960 30000 6 trzf2_clk
port 374 nsew signal output
rlabel metal2 s 71232 29600 71288 30000 6 trzf2_ena
port 375 nsew signal output
rlabel metal2 s 116928 29600 116984 30000 6 trzf2_io_in[0]
port 376 nsew signal output
rlabel metal2 s 110208 29600 110264 30000 6 trzf2_io_in[10]
port 377 nsew signal output
rlabel metal2 s 109536 29600 109592 30000 6 trzf2_io_in[11]
port 378 nsew signal output
rlabel metal2 s 108864 29600 108920 30000 6 trzf2_io_in[12]
port 379 nsew signal output
rlabel metal2 s 108192 29600 108248 30000 6 trzf2_io_in[13]
port 380 nsew signal output
rlabel metal2 s 107520 29600 107576 30000 6 trzf2_io_in[14]
port 381 nsew signal output
rlabel metal2 s 106848 29600 106904 30000 6 trzf2_io_in[15]
port 382 nsew signal output
rlabel metal2 s 106176 29600 106232 30000 6 trzf2_io_in[16]
port 383 nsew signal output
rlabel metal2 s 105504 29600 105560 30000 6 trzf2_io_in[17]
port 384 nsew signal output
rlabel metal2 s 104832 29600 104888 30000 6 trzf2_io_in[18]
port 385 nsew signal output
rlabel metal2 s 104160 29600 104216 30000 6 trzf2_io_in[19]
port 386 nsew signal output
rlabel metal2 s 116256 29600 116312 30000 6 trzf2_io_in[1]
port 387 nsew signal output
rlabel metal2 s 103488 29600 103544 30000 6 trzf2_io_in[20]
port 388 nsew signal output
rlabel metal2 s 102816 29600 102872 30000 6 trzf2_io_in[21]
port 389 nsew signal output
rlabel metal2 s 102144 29600 102200 30000 6 trzf2_io_in[22]
port 390 nsew signal output
rlabel metal2 s 101472 29600 101528 30000 6 trzf2_io_in[23]
port 391 nsew signal output
rlabel metal2 s 100800 29600 100856 30000 6 trzf2_io_in[24]
port 392 nsew signal output
rlabel metal2 s 100128 29600 100184 30000 6 trzf2_io_in[25]
port 393 nsew signal output
rlabel metal2 s 99456 29600 99512 30000 6 trzf2_io_in[26]
port 394 nsew signal output
rlabel metal2 s 98784 29600 98840 30000 6 trzf2_io_in[27]
port 395 nsew signal output
rlabel metal2 s 98112 29600 98168 30000 6 trzf2_io_in[28]
port 396 nsew signal output
rlabel metal2 s 97440 29600 97496 30000 6 trzf2_io_in[29]
port 397 nsew signal output
rlabel metal2 s 115584 29600 115640 30000 6 trzf2_io_in[2]
port 398 nsew signal output
rlabel metal2 s 96768 29600 96824 30000 6 trzf2_io_in[30]
port 399 nsew signal output
rlabel metal2 s 96096 29600 96152 30000 6 trzf2_io_in[31]
port 400 nsew signal output
rlabel metal2 s 95424 29600 95480 30000 6 trzf2_io_in[32]
port 401 nsew signal output
rlabel metal2 s 94752 29600 94808 30000 6 trzf2_io_in[33]
port 402 nsew signal output
rlabel metal2 s 94080 29600 94136 30000 6 trzf2_io_in[34]
port 403 nsew signal output
rlabel metal2 s 93408 29600 93464 30000 6 trzf2_io_in[35]
port 404 nsew signal output
rlabel metal2 s 92736 29600 92792 30000 6 trzf2_io_in[36]
port 405 nsew signal output
rlabel metal2 s 92064 29600 92120 30000 6 trzf2_io_in[37]
port 406 nsew signal output
rlabel metal2 s 114912 29600 114968 30000 6 trzf2_io_in[3]
port 407 nsew signal output
rlabel metal2 s 114240 29600 114296 30000 6 trzf2_io_in[4]
port 408 nsew signal output
rlabel metal2 s 113568 29600 113624 30000 6 trzf2_io_in[5]
port 409 nsew signal output
rlabel metal2 s 112896 29600 112952 30000 6 trzf2_io_in[6]
port 410 nsew signal output
rlabel metal2 s 112224 29600 112280 30000 6 trzf2_io_in[7]
port 411 nsew signal output
rlabel metal2 s 111552 29600 111608 30000 6 trzf2_io_in[8]
port 412 nsew signal output
rlabel metal2 s 110880 29600 110936 30000 6 trzf2_io_in[9]
port 413 nsew signal output
rlabel metal2 s 81312 29600 81368 30000 6 trzf2_la_in[0]
port 414 nsew signal output
rlabel metal2 s 74592 29600 74648 30000 6 trzf2_la_in[10]
port 415 nsew signal output
rlabel metal2 s 73920 29600 73976 30000 6 trzf2_la_in[11]
port 416 nsew signal output
rlabel metal2 s 73248 29600 73304 30000 6 trzf2_la_in[12]
port 417 nsew signal output
rlabel metal2 s 80640 29600 80696 30000 6 trzf2_la_in[1]
port 418 nsew signal output
rlabel metal2 s 79968 29600 80024 30000 6 trzf2_la_in[2]
port 419 nsew signal output
rlabel metal2 s 79296 29600 79352 30000 6 trzf2_la_in[3]
port 420 nsew signal output
rlabel metal2 s 78624 29600 78680 30000 6 trzf2_la_in[4]
port 421 nsew signal output
rlabel metal2 s 77952 29600 78008 30000 6 trzf2_la_in[5]
port 422 nsew signal output
rlabel metal2 s 77280 29600 77336 30000 6 trzf2_la_in[6]
port 423 nsew signal output
rlabel metal2 s 76608 29600 76664 30000 6 trzf2_la_in[7]
port 424 nsew signal output
rlabel metal2 s 75936 29600 75992 30000 6 trzf2_la_in[8]
port 425 nsew signal output
rlabel metal2 s 75264 29600 75320 30000 6 trzf2_la_in[9]
port 426 nsew signal output
rlabel metal2 s 83328 29600 83384 30000 6 trzf2_o_gpout[0]
port 427 nsew signal input
rlabel metal2 s 82656 29600 82712 30000 6 trzf2_o_gpout[1]
port 428 nsew signal input
rlabel metal2 s 81984 29600 82040 30000 6 trzf2_o_gpout[2]
port 429 nsew signal input
rlabel metal2 s 91392 29600 91448 30000 6 trzf2_o_hsync
port 430 nsew signal input
rlabel metal2 s 90048 29600 90104 30000 6 trzf2_o_rgb[0]
port 431 nsew signal input
rlabel metal2 s 89376 29600 89432 30000 6 trzf2_o_rgb[1]
port 432 nsew signal input
rlabel metal2 s 88704 29600 88760 30000 6 trzf2_o_rgb[2]
port 433 nsew signal input
rlabel metal2 s 88032 29600 88088 30000 6 trzf2_o_rgb[3]
port 434 nsew signal input
rlabel metal2 s 87360 29600 87416 30000 6 trzf2_o_rgb[4]
port 435 nsew signal input
rlabel metal2 s 86688 29600 86744 30000 6 trzf2_o_rgb[5]
port 436 nsew signal input
rlabel metal2 s 86016 29600 86072 30000 6 trzf2_o_tex_csb
port 437 nsew signal input
rlabel metal2 s 84000 29600 84056 30000 6 trzf2_o_tex_oeb0
port 438 nsew signal input
rlabel metal2 s 84672 29600 84728 30000 6 trzf2_o_tex_out0
port 439 nsew signal input
rlabel metal2 s 85344 29600 85400 30000 6 trzf2_o_tex_sclk
port 440 nsew signal input
rlabel metal2 s 90720 29600 90776 30000 6 trzf2_o_vsync
port 441 nsew signal input
rlabel metal2 s 72576 29600 72632 30000 6 trzf2_rst
port 442 nsew signal output
rlabel metal2 s 4032 29600 4088 30000 6 trzf_clk
port 443 nsew signal output
rlabel metal2 s 3360 29600 3416 30000 6 trzf_ena
port 444 nsew signal output
rlabel metal2 s 49056 29600 49112 30000 6 trzf_io_in[0]
port 445 nsew signal output
rlabel metal2 s 42336 29600 42392 30000 6 trzf_io_in[10]
port 446 nsew signal output
rlabel metal2 s 41664 29600 41720 30000 6 trzf_io_in[11]
port 447 nsew signal output
rlabel metal2 s 40992 29600 41048 30000 6 trzf_io_in[12]
port 448 nsew signal output
rlabel metal2 s 40320 29600 40376 30000 6 trzf_io_in[13]
port 449 nsew signal output
rlabel metal2 s 39648 29600 39704 30000 6 trzf_io_in[14]
port 450 nsew signal output
rlabel metal2 s 38976 29600 39032 30000 6 trzf_io_in[15]
port 451 nsew signal output
rlabel metal2 s 38304 29600 38360 30000 6 trzf_io_in[16]
port 452 nsew signal output
rlabel metal2 s 37632 29600 37688 30000 6 trzf_io_in[17]
port 453 nsew signal output
rlabel metal2 s 36960 29600 37016 30000 6 trzf_io_in[18]
port 454 nsew signal output
rlabel metal2 s 36288 29600 36344 30000 6 trzf_io_in[19]
port 455 nsew signal output
rlabel metal2 s 48384 29600 48440 30000 6 trzf_io_in[1]
port 456 nsew signal output
rlabel metal2 s 35616 29600 35672 30000 6 trzf_io_in[20]
port 457 nsew signal output
rlabel metal2 s 34944 29600 35000 30000 6 trzf_io_in[21]
port 458 nsew signal output
rlabel metal2 s 34272 29600 34328 30000 6 trzf_io_in[22]
port 459 nsew signal output
rlabel metal2 s 33600 29600 33656 30000 6 trzf_io_in[23]
port 460 nsew signal output
rlabel metal2 s 32928 29600 32984 30000 6 trzf_io_in[24]
port 461 nsew signal output
rlabel metal2 s 32256 29600 32312 30000 6 trzf_io_in[25]
port 462 nsew signal output
rlabel metal2 s 31584 29600 31640 30000 6 trzf_io_in[26]
port 463 nsew signal output
rlabel metal2 s 30912 29600 30968 30000 6 trzf_io_in[27]
port 464 nsew signal output
rlabel metal2 s 30240 29600 30296 30000 6 trzf_io_in[28]
port 465 nsew signal output
rlabel metal2 s 29568 29600 29624 30000 6 trzf_io_in[29]
port 466 nsew signal output
rlabel metal2 s 47712 29600 47768 30000 6 trzf_io_in[2]
port 467 nsew signal output
rlabel metal2 s 28896 29600 28952 30000 6 trzf_io_in[30]
port 468 nsew signal output
rlabel metal2 s 28224 29600 28280 30000 6 trzf_io_in[31]
port 469 nsew signal output
rlabel metal2 s 27552 29600 27608 30000 6 trzf_io_in[32]
port 470 nsew signal output
rlabel metal2 s 26880 29600 26936 30000 6 trzf_io_in[33]
port 471 nsew signal output
rlabel metal2 s 26208 29600 26264 30000 6 trzf_io_in[34]
port 472 nsew signal output
rlabel metal2 s 25536 29600 25592 30000 6 trzf_io_in[35]
port 473 nsew signal output
rlabel metal2 s 24864 29600 24920 30000 6 trzf_io_in[36]
port 474 nsew signal output
rlabel metal2 s 24192 29600 24248 30000 6 trzf_io_in[37]
port 475 nsew signal output
rlabel metal2 s 47040 29600 47096 30000 6 trzf_io_in[3]
port 476 nsew signal output
rlabel metal2 s 46368 29600 46424 30000 6 trzf_io_in[4]
port 477 nsew signal output
rlabel metal2 s 45696 29600 45752 30000 6 trzf_io_in[5]
port 478 nsew signal output
rlabel metal2 s 45024 29600 45080 30000 6 trzf_io_in[6]
port 479 nsew signal output
rlabel metal2 s 44352 29600 44408 30000 6 trzf_io_in[7]
port 480 nsew signal output
rlabel metal2 s 43680 29600 43736 30000 6 trzf_io_in[8]
port 481 nsew signal output
rlabel metal2 s 43008 29600 43064 30000 6 trzf_io_in[9]
port 482 nsew signal output
rlabel metal2 s 13440 29600 13496 30000 6 trzf_la_in[0]
port 483 nsew signal output
rlabel metal2 s 6720 29600 6776 30000 6 trzf_la_in[10]
port 484 nsew signal output
rlabel metal2 s 6048 29600 6104 30000 6 trzf_la_in[11]
port 485 nsew signal output
rlabel metal2 s 5376 29600 5432 30000 6 trzf_la_in[12]
port 486 nsew signal output
rlabel metal2 s 12768 29600 12824 30000 6 trzf_la_in[1]
port 487 nsew signal output
rlabel metal2 s 12096 29600 12152 30000 6 trzf_la_in[2]
port 488 nsew signal output
rlabel metal2 s 11424 29600 11480 30000 6 trzf_la_in[3]
port 489 nsew signal output
rlabel metal2 s 10752 29600 10808 30000 6 trzf_la_in[4]
port 490 nsew signal output
rlabel metal2 s 10080 29600 10136 30000 6 trzf_la_in[5]
port 491 nsew signal output
rlabel metal2 s 9408 29600 9464 30000 6 trzf_la_in[6]
port 492 nsew signal output
rlabel metal2 s 8736 29600 8792 30000 6 trzf_la_in[7]
port 493 nsew signal output
rlabel metal2 s 8064 29600 8120 30000 6 trzf_la_in[8]
port 494 nsew signal output
rlabel metal2 s 7392 29600 7448 30000 6 trzf_la_in[9]
port 495 nsew signal output
rlabel metal2 s 15456 29600 15512 30000 6 trzf_o_gpout[0]
port 496 nsew signal input
rlabel metal2 s 14784 29600 14840 30000 6 trzf_o_gpout[1]
port 497 nsew signal input
rlabel metal2 s 14112 29600 14168 30000 6 trzf_o_gpout[2]
port 498 nsew signal input
rlabel metal2 s 23520 29600 23576 30000 6 trzf_o_hsync
port 499 nsew signal input
rlabel metal2 s 22176 29600 22232 30000 6 trzf_o_rgb[0]
port 500 nsew signal input
rlabel metal2 s 21504 29600 21560 30000 6 trzf_o_rgb[1]
port 501 nsew signal input
rlabel metal2 s 20832 29600 20888 30000 6 trzf_o_rgb[2]
port 502 nsew signal input
rlabel metal2 s 20160 29600 20216 30000 6 trzf_o_rgb[3]
port 503 nsew signal input
rlabel metal2 s 19488 29600 19544 30000 6 trzf_o_rgb[4]
port 504 nsew signal input
rlabel metal2 s 18816 29600 18872 30000 6 trzf_o_rgb[5]
port 505 nsew signal input
rlabel metal2 s 18144 29600 18200 30000 6 trzf_o_tex_csb
port 506 nsew signal input
rlabel metal2 s 16128 29600 16184 30000 6 trzf_o_tex_oeb0
port 507 nsew signal input
rlabel metal2 s 16800 29600 16856 30000 6 trzf_o_tex_out0
port 508 nsew signal input
rlabel metal2 s 17472 29600 17528 30000 6 trzf_o_tex_sclk
port 509 nsew signal input
rlabel metal2 s 22848 29600 22904 30000 6 trzf_o_vsync
port 510 nsew signal input
rlabel metal2 s 4704 29600 4760 30000 6 trzf_rst
port 511 nsew signal output
rlabel metal2 s 52752 0 52808 400 6 uri_clk
port 512 nsew signal output
rlabel metal2 s 54096 0 54152 400 6 uri_ena
port 513 nsew signal output
rlabel metal2 s 54768 0 54824 400 6 uri_io_in[0]
port 514 nsew signal output
rlabel metal2 s 74928 0 74984 400 6 uri_io_in[10]
port 515 nsew signal output
rlabel metal2 s 76944 0 77000 400 6 uri_io_in[11]
port 516 nsew signal output
rlabel metal2 s 78960 0 79016 400 6 uri_io_in[12]
port 517 nsew signal output
rlabel metal2 s 80976 0 81032 400 6 uri_io_in[13]
port 518 nsew signal output
rlabel metal2 s 82992 0 83048 400 6 uri_io_in[14]
port 519 nsew signal output
rlabel metal2 s 85008 0 85064 400 6 uri_io_in[15]
port 520 nsew signal output
rlabel metal2 s 87024 0 87080 400 6 uri_io_in[16]
port 521 nsew signal output
rlabel metal2 s 89040 0 89096 400 6 uri_io_in[17]
port 522 nsew signal output
rlabel metal2 s 91056 0 91112 400 6 uri_io_in[18]
port 523 nsew signal output
rlabel metal2 s 93072 0 93128 400 6 uri_io_in[19]
port 524 nsew signal output
rlabel metal2 s 56784 0 56840 400 6 uri_io_in[1]
port 525 nsew signal output
rlabel metal2 s 93744 0 93800 400 6 uri_io_in[20]
port 526 nsew signal output
rlabel metal2 s 94416 0 94472 400 6 uri_io_in[21]
port 527 nsew signal output
rlabel metal2 s 95088 0 95144 400 6 uri_io_in[22]
port 528 nsew signal output
rlabel metal2 s 95760 0 95816 400 6 uri_io_in[23]
port 529 nsew signal output
rlabel metal2 s 96432 0 96488 400 6 uri_io_in[24]
port 530 nsew signal output
rlabel metal2 s 97104 0 97160 400 6 uri_io_in[25]
port 531 nsew signal output
rlabel metal2 s 97776 0 97832 400 6 uri_io_in[26]
port 532 nsew signal output
rlabel metal2 s 98448 0 98504 400 6 uri_io_in[27]
port 533 nsew signal output
rlabel metal2 s 99120 0 99176 400 6 uri_io_in[28]
port 534 nsew signal output
rlabel metal2 s 99792 0 99848 400 6 uri_io_in[29]
port 535 nsew signal output
rlabel metal2 s 58800 0 58856 400 6 uri_io_in[2]
port 536 nsew signal output
rlabel metal2 s 100464 0 100520 400 6 uri_io_in[30]
port 537 nsew signal output
rlabel metal2 s 101136 0 101192 400 6 uri_io_in[31]
port 538 nsew signal output
rlabel metal2 s 101808 0 101864 400 6 uri_io_in[32]
port 539 nsew signal output
rlabel metal2 s 102480 0 102536 400 6 uri_io_in[33]
port 540 nsew signal output
rlabel metal2 s 103152 0 103208 400 6 uri_io_in[34]
port 541 nsew signal output
rlabel metal2 s 103824 0 103880 400 6 uri_io_in[35]
port 542 nsew signal output
rlabel metal2 s 104496 0 104552 400 6 uri_io_in[36]
port 543 nsew signal output
rlabel metal2 s 105168 0 105224 400 6 uri_io_in[37]
port 544 nsew signal output
rlabel metal2 s 60816 0 60872 400 6 uri_io_in[3]
port 545 nsew signal output
rlabel metal2 s 62832 0 62888 400 6 uri_io_in[4]
port 546 nsew signal output
rlabel metal2 s 64848 0 64904 400 6 uri_io_in[5]
port 547 nsew signal output
rlabel metal2 s 66864 0 66920 400 6 uri_io_in[6]
port 548 nsew signal output
rlabel metal2 s 68880 0 68936 400 6 uri_io_in[7]
port 549 nsew signal output
rlabel metal2 s 70896 0 70952 400 6 uri_io_in[8]
port 550 nsew signal output
rlabel metal2 s 72912 0 72968 400 6 uri_io_in[9]
port 551 nsew signal output
rlabel metal2 s 55440 0 55496 400 6 uri_io_oeb[0]
port 552 nsew signal input
rlabel metal2 s 75600 0 75656 400 6 uri_io_oeb[10]
port 553 nsew signal input
rlabel metal2 s 77616 0 77672 400 6 uri_io_oeb[11]
port 554 nsew signal input
rlabel metal2 s 79632 0 79688 400 6 uri_io_oeb[12]
port 555 nsew signal input
rlabel metal2 s 81648 0 81704 400 6 uri_io_oeb[13]
port 556 nsew signal input
rlabel metal2 s 83664 0 83720 400 6 uri_io_oeb[14]
port 557 nsew signal input
rlabel metal2 s 85680 0 85736 400 6 uri_io_oeb[15]
port 558 nsew signal input
rlabel metal2 s 87696 0 87752 400 6 uri_io_oeb[16]
port 559 nsew signal input
rlabel metal2 s 89712 0 89768 400 6 uri_io_oeb[17]
port 560 nsew signal input
rlabel metal2 s 91728 0 91784 400 6 uri_io_oeb[18]
port 561 nsew signal input
rlabel metal2 s 57456 0 57512 400 6 uri_io_oeb[1]
port 562 nsew signal input
rlabel metal2 s 59472 0 59528 400 6 uri_io_oeb[2]
port 563 nsew signal input
rlabel metal2 s 61488 0 61544 400 6 uri_io_oeb[3]
port 564 nsew signal input
rlabel metal2 s 63504 0 63560 400 6 uri_io_oeb[4]
port 565 nsew signal input
rlabel metal2 s 65520 0 65576 400 6 uri_io_oeb[5]
port 566 nsew signal input
rlabel metal2 s 67536 0 67592 400 6 uri_io_oeb[6]
port 567 nsew signal input
rlabel metal2 s 69552 0 69608 400 6 uri_io_oeb[7]
port 568 nsew signal input
rlabel metal2 s 71568 0 71624 400 6 uri_io_oeb[8]
port 569 nsew signal input
rlabel metal2 s 73584 0 73640 400 6 uri_io_oeb[9]
port 570 nsew signal input
rlabel metal2 s 56112 0 56168 400 6 uri_io_out[0]
port 571 nsew signal input
rlabel metal2 s 76272 0 76328 400 6 uri_io_out[10]
port 572 nsew signal input
rlabel metal2 s 78288 0 78344 400 6 uri_io_out[11]
port 573 nsew signal input
rlabel metal2 s 80304 0 80360 400 6 uri_io_out[12]
port 574 nsew signal input
rlabel metal2 s 82320 0 82376 400 6 uri_io_out[13]
port 575 nsew signal input
rlabel metal2 s 84336 0 84392 400 6 uri_io_out[14]
port 576 nsew signal input
rlabel metal2 s 86352 0 86408 400 6 uri_io_out[15]
port 577 nsew signal input
rlabel metal2 s 88368 0 88424 400 6 uri_io_out[16]
port 578 nsew signal input
rlabel metal2 s 90384 0 90440 400 6 uri_io_out[17]
port 579 nsew signal input
rlabel metal2 s 92400 0 92456 400 6 uri_io_out[18]
port 580 nsew signal input
rlabel metal2 s 58128 0 58184 400 6 uri_io_out[1]
port 581 nsew signal input
rlabel metal2 s 60144 0 60200 400 6 uri_io_out[2]
port 582 nsew signal input
rlabel metal2 s 62160 0 62216 400 6 uri_io_out[3]
port 583 nsew signal input
rlabel metal2 s 64176 0 64232 400 6 uri_io_out[4]
port 584 nsew signal input
rlabel metal2 s 66192 0 66248 400 6 uri_io_out[5]
port 585 nsew signal input
rlabel metal2 s 68208 0 68264 400 6 uri_io_out[6]
port 586 nsew signal input
rlabel metal2 s 70224 0 70280 400 6 uri_io_out[7]
port 587 nsew signal input
rlabel metal2 s 72240 0 72296 400 6 uri_io_out[8]
port 588 nsew signal input
rlabel metal2 s 74256 0 74312 400 6 uri_io_out[9]
port 589 nsew signal input
rlabel metal2 s 53424 0 53480 400 6 uri_rst
port 590 nsew signal output
rlabel metal4 s 2224 1538 2384 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 28254 6 vdd
port 591 nsew power bidirectional
rlabel metal2 s 144480 29600 144536 30000 6 vgasp_clk
port 592 nsew signal output
rlabel metal2 s 170688 29600 170744 30000 6 vgasp_io_in[0]
port 593 nsew signal output
rlabel metal2 s 163968 29600 164024 30000 6 vgasp_io_in[10]
port 594 nsew signal output
rlabel metal2 s 163296 29600 163352 30000 6 vgasp_io_in[11]
port 595 nsew signal output
rlabel metal2 s 162624 29600 162680 30000 6 vgasp_io_in[12]
port 596 nsew signal output
rlabel metal2 s 161952 29600 162008 30000 6 vgasp_io_in[13]
port 597 nsew signal output
rlabel metal2 s 161280 29600 161336 30000 6 vgasp_io_in[14]
port 598 nsew signal output
rlabel metal2 s 160608 29600 160664 30000 6 vgasp_io_in[15]
port 599 nsew signal output
rlabel metal2 s 159936 29600 159992 30000 6 vgasp_io_in[16]
port 600 nsew signal output
rlabel metal2 s 159264 29600 159320 30000 6 vgasp_io_in[17]
port 601 nsew signal output
rlabel metal2 s 158592 29600 158648 30000 6 vgasp_io_in[18]
port 602 nsew signal output
rlabel metal2 s 157920 29600 157976 30000 6 vgasp_io_in[19]
port 603 nsew signal output
rlabel metal2 s 170016 29600 170072 30000 6 vgasp_io_in[1]
port 604 nsew signal output
rlabel metal2 s 157248 29600 157304 30000 6 vgasp_io_in[20]
port 605 nsew signal output
rlabel metal2 s 156576 29600 156632 30000 6 vgasp_io_in[21]
port 606 nsew signal output
rlabel metal2 s 155904 29600 155960 30000 6 vgasp_io_in[22]
port 607 nsew signal output
rlabel metal2 s 155232 29600 155288 30000 6 vgasp_io_in[23]
port 608 nsew signal output
rlabel metal2 s 154560 29600 154616 30000 6 vgasp_io_in[24]
port 609 nsew signal output
rlabel metal2 s 153888 29600 153944 30000 6 vgasp_io_in[25]
port 610 nsew signal output
rlabel metal2 s 153216 29600 153272 30000 6 vgasp_io_in[26]
port 611 nsew signal output
rlabel metal2 s 152544 29600 152600 30000 6 vgasp_io_in[27]
port 612 nsew signal output
rlabel metal2 s 151872 29600 151928 30000 6 vgasp_io_in[28]
port 613 nsew signal output
rlabel metal2 s 151200 29600 151256 30000 6 vgasp_io_in[29]
port 614 nsew signal output
rlabel metal2 s 169344 29600 169400 30000 6 vgasp_io_in[2]
port 615 nsew signal output
rlabel metal2 s 150528 29600 150584 30000 6 vgasp_io_in[30]
port 616 nsew signal output
rlabel metal2 s 149856 29600 149912 30000 6 vgasp_io_in[31]
port 617 nsew signal output
rlabel metal2 s 149184 29600 149240 30000 6 vgasp_io_in[32]
port 618 nsew signal output
rlabel metal2 s 148512 29600 148568 30000 6 vgasp_io_in[33]
port 619 nsew signal output
rlabel metal2 s 147840 29600 147896 30000 6 vgasp_io_in[34]
port 620 nsew signal output
rlabel metal2 s 147168 29600 147224 30000 6 vgasp_io_in[35]
port 621 nsew signal output
rlabel metal2 s 146496 29600 146552 30000 6 vgasp_io_in[36]
port 622 nsew signal output
rlabel metal2 s 145824 29600 145880 30000 6 vgasp_io_in[37]
port 623 nsew signal output
rlabel metal2 s 168672 29600 168728 30000 6 vgasp_io_in[3]
port 624 nsew signal output
rlabel metal2 s 168000 29600 168056 30000 6 vgasp_io_in[4]
port 625 nsew signal output
rlabel metal2 s 167328 29600 167384 30000 6 vgasp_io_in[5]
port 626 nsew signal output
rlabel metal2 s 166656 29600 166712 30000 6 vgasp_io_in[6]
port 627 nsew signal output
rlabel metal2 s 165984 29600 166040 30000 6 vgasp_io_in[7]
port 628 nsew signal output
rlabel metal2 s 165312 29600 165368 30000 6 vgasp_io_in[8]
port 629 nsew signal output
rlabel metal2 s 164640 29600 164696 30000 6 vgasp_io_in[9]
port 630 nsew signal output
rlabel metal2 s 145152 29600 145208 30000 6 vgasp_rst
port 631 nsew signal output
rlabel metal2 s 186816 29600 186872 30000 6 vgasp_uio_oe[0]
port 632 nsew signal input
rlabel metal2 s 186144 29600 186200 30000 6 vgasp_uio_oe[1]
port 633 nsew signal input
rlabel metal2 s 185472 29600 185528 30000 6 vgasp_uio_oe[2]
port 634 nsew signal input
rlabel metal2 s 184800 29600 184856 30000 6 vgasp_uio_oe[3]
port 635 nsew signal input
rlabel metal2 s 184128 29600 184184 30000 6 vgasp_uio_oe[4]
port 636 nsew signal input
rlabel metal2 s 183456 29600 183512 30000 6 vgasp_uio_oe[5]
port 637 nsew signal input
rlabel metal2 s 182784 29600 182840 30000 6 vgasp_uio_oe[6]
port 638 nsew signal input
rlabel metal2 s 182112 29600 182168 30000 6 vgasp_uio_oe[7]
port 639 nsew signal input
rlabel metal2 s 181440 29600 181496 30000 6 vgasp_uio_out[0]
port 640 nsew signal input
rlabel metal2 s 180768 29600 180824 30000 6 vgasp_uio_out[1]
port 641 nsew signal input
rlabel metal2 s 180096 29600 180152 30000 6 vgasp_uio_out[2]
port 642 nsew signal input
rlabel metal2 s 179424 29600 179480 30000 6 vgasp_uio_out[3]
port 643 nsew signal input
rlabel metal2 s 178752 29600 178808 30000 6 vgasp_uio_out[4]
port 644 nsew signal input
rlabel metal2 s 178080 29600 178136 30000 6 vgasp_uio_out[5]
port 645 nsew signal input
rlabel metal2 s 177408 29600 177464 30000 6 vgasp_uio_out[6]
port 646 nsew signal input
rlabel metal2 s 176736 29600 176792 30000 6 vgasp_uio_out[7]
port 647 nsew signal input
rlabel metal2 s 176064 29600 176120 30000 6 vgasp_uo_out[0]
port 648 nsew signal input
rlabel metal2 s 175392 29600 175448 30000 6 vgasp_uo_out[1]
port 649 nsew signal input
rlabel metal2 s 174720 29600 174776 30000 6 vgasp_uo_out[2]
port 650 nsew signal input
rlabel metal2 s 174048 29600 174104 30000 6 vgasp_uo_out[3]
port 651 nsew signal input
rlabel metal2 s 173376 29600 173432 30000 6 vgasp_uo_out[4]
port 652 nsew signal input
rlabel metal2 s 172704 29600 172760 30000 6 vgasp_uo_out[5]
port 653 nsew signal input
rlabel metal2 s 172032 29600 172088 30000 6 vgasp_uo_out[6]
port 654 nsew signal input
rlabel metal2 s 171360 29600 171416 30000 6 vgasp_uo_out[7]
port 655 nsew signal input
rlabel metal4 s 9904 1538 10064 28254 6 vss
port 656 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 28254 6 vss
port 656 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 28254 6 vss
port 656 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 28254 6 vss
port 656 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 28254 6 vss
port 656 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 28254 6 vss
port 656 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 28254 6 vss
port 656 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 28254 6 vss
port 656 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 28254 6 vss
port 656 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 28254 6 vss
port 656 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 28254 6 vss
port 656 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 28254 6 vss
port 656 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 28254 6 vss
port 656 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 28254 6 vss
port 656 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 28254 6 vss
port 656 nsew ground bidirectional
rlabel metal3 s 0 2576 400 2632 6 wb_clk_i
port 657 nsew signal input
rlabel metal3 s 0 2016 400 2072 6 wb_rst_i
port 658 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 240000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4664662
string GDS_FILE /home/zerotoasic/anton/algofoogle-multi-caravel/openlane/top_design_mux/runs/23_12_12_00_07/results/signoff/top_design_mux.magic.gds
string GDS_START 299144
<< end >>

